
package picorv32_pkg;

  parameter CPU_CLK   = 50_000_000;   //Default CPU frequency on FPGA
  parameter SRAM_BAUD_RATE = 9600;          //Default Baud rate for programming on the run via UART

  parameter [ 0:0] ENABLE_COUNTERS = 1            ;
  parameter [ 0:0] ENABLE_COUNTERS64 = 0          ;
  parameter [ 0:0] ENABLE_REGS_16_31 = 1          ;
  parameter [ 0:0] ENABLE_REGS_DUALPORT = 1       ;
  parameter [ 0:0] LATCHED_MEM_RDATA = 0          ;
  parameter [ 0:0] TWO_STAGE_SHIFT = 1            ;
  parameter [ 0:0] BARREL_SHIFTER = 0             ;
  parameter [ 0:0] TWO_CYCLE_COMPARE = 0          ;
  parameter [ 0:0] TWO_CYCLE_ALU = 0              ;
  parameter [ 0:0] COMPRESSED_ISA = 1             ;
  parameter [ 0:0] CATCH_MISALIGN = 1             ;
  parameter [ 0:0] CATCH_ILLINSN = 1              ;
  parameter [ 0:0] ENABLE_PCPI = 0                ;
  parameter [ 0:0] ENABLE_MUL = 1                 ;
  parameter [ 0:0] ENABLE_FAST_MUL = 0            ;
  parameter [ 0:0] ENABLE_DIV = 1                 ;
  parameter [ 0:0] ENABLE_IRQ = 1                 ;
  parameter [ 0:0] ENABLE_IRQ_QREGS = 0           ;
  parameter [ 0:0] ENABLE_IRQ_TIMER = 0           ;
  parameter [ 0:0] ENABLE_TRACE = 0               ;
  parameter [ 0:0] REGS_INIT_ZERO = 0             ;
  parameter [31:0] MASKED_IRQ = 32'h 0000_0000    ;
  parameter [31:0] LATCHED_IRQ = 32'h ffff_ffff   ;

  //parameter BOOT_FILE = ""; // /home/yunus.eryilmaz/sim_workspace/picosoc/sw/outputs/hex/picosoc_test.hex
  parameter integer RAM_DEPTH = 131072;
   
  parameter [31:0] PROGADDR_RESET = 32'h4000_0000; // RAM base addr
  parameter [31:0] STACKADDR = PROGADDR_RESET + (4*RAM_DEPTH);       // end of memory
  parameter [31:0] PROGADDR_IRQ      = 32'h0000_0000;
  parameter [31:0] UART_BASE_ADDR    = 32'h2000_0000;
  parameter [31:0] UART_MASK_ADDR    = 32'h0000_000f;
  parameter [31:0] SPI_BASE_ADDR     = 32'h2001_0000;
  parameter [31:0] SPI_MASK_ADDR     = 32'h0000_00ff;
  parameter [31:0] PWM_BASE_ADDR     = 32'h2002_0000;
  parameter [31:0] PWM_MASK_ADDR     = 32'h0000_00ff;
  parameter [31:0] TIMER_BASE_ADDR   = 32'h2003_0000;
  parameter [31:0] TIMER_MASK_ADDR   = 32'h0000_000f;
  parameter [31:0] I2C_BASE_ADDR     = 32'h2004_0000;
  parameter [31:0] I2C_MASK_ADDR     = 32'h0000_00ff;
  parameter [31:0] SRAM_BASE_ADDR    = 32'h4000_0000;
  parameter [31:0] SRAM_MASK_ADDR    = 32'h000f_ffff;
  parameter [31:0] EFPGA_BASE_ADDR   = 32'h4200_0000;
  parameter [31:0] EFPGA_MASK_ADDR   = 32'h000f_ffff;

  parameter [31:0] CHIP_IO_BASE_ADDR = SPI_BASE_ADDR + SPI_MASK_ADDR;
  parameter [31:0] CHIP_IO_MASK_ADDR = SRAM_BASE_ADDR + SRAM_MASK_ADDR;
   
  typedef struct packed {
    logic [31:0] a_adr;
    logic [31:0] a_dat;
    logic        a_we ;
    logic [ 3:0] a_sel;
    logic        a_stb;
    logic        a_cyc;    
  } wb_h2d_t;
 
  typedef struct packed {
    logic [31:0] d_dat;
    logic        d_ack;    
  } wb_d2h_t;

  
endpackage
