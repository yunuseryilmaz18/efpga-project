`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.06.2022 10:48:02
// Design Name: 
// Module Name: picosoc_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module picosoc_tb();

reg clk_in1;
reg rst_ni;

wire uart_tx_o;
reg  uart_rx_i;

reg  sram_rx_i;
wire sram_prog_led_o;

wire cio_sck_o ;
wire cio_csb_o ;
wire cio_mosi_o ;
wire cio_miso_i ;

parameter BOOT_FILE = "/home/yunus.eryilmaz/sim_workspace/picosoc/sw/outputs/hex/picosoc_system_efpga.hex";

picosoc #(.BOOT_FILE(BOOT_FILE))
	uut (
	.clk_in1,
	.rst_ni,

	.uart_tx_o,
	.uart_rx_i,
	
	.sram_rx_i,           
	.sram_prog_led_o,
	   
    .cio_sck_o ,
    .cio_csb_o ,
    .cio_mosi_o,
    .cio_miso_i
);

wire   WPn  ;
wire   HOLDn;
assign WPn   = 1'b1;
assign HOLDn = 1'b1;

initial begin
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_1__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = 64'b1111111100000000111111110000000000000000000000000000000000000000;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = 64'b0000000011111111000000001111111111111111111111111111111111111111;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b010;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b101;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0010000000100000;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1101111111011111;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0010000001000000;
	force uut.u_efpga.FPGA.grid_clb_2__1_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1101111110111111;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_8.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_out[0:63] = {64{1'b0}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.logical_tile_clb_mode_default__fle_mode_physical__ble6_mode_default__lut6_0.lut6_DFFR_mem.mem_outb[0:63] = {64{1'b1}};
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_out[0:2] = 3'b001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_9.logical_tile_clb_mode_default__fle_mode_physical__ble6_0.mem_ble6_out_0.mem_outb[0:2] = 3'b110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_4_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_5_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_6_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_7_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_8_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_0.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_1.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_2.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_3.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_4.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_out[0:15] = 16'b0000000000000001;
	force uut.u_efpga.FPGA.grid_clb_2__2_.logical_tile_clb_mode_clb__0.mem_fle_9_in_5.mem_outb[0:15] = 16'b1111111111111110;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_1__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_top_2__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_right_3__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_out[0] = 1'b1;
	force uut.u_efpga.FPGA.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFFR_mem.mem_outb[0] = 1'b0;
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__1_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_0__1_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_0__1_.mem_top_track_8.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_0__1_.mem_top_track_8.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_0__1_.mem_right_track_2.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_0__1_.mem_right_track_2.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_0__1_.mem_right_track_4.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_0__1_.mem_right_track_4.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_0__1_.mem_right_track_6.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_0__1_.mem_right_track_6.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_0__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00100100;
	force uut.u_efpga.FPGA.sb_0__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11011011;
	force uut.u_efpga.FPGA.sb_0__1_.mem_bottom_track_9.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_0__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_0.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_0.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_0__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_0.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_0.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_8.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_1__0_.mem_top_track_8.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_1__0_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__0_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__0_.mem_right_track_8.mem_out[0:7] = 8'b10001000;
	force uut.u_efpga.FPGA.sb_1__0_.mem_right_track_8.mem_outb[0:7] = 8'b01110111;
	force uut.u_efpga.FPGA.sb_1__0_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__0_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__0_.mem_left_track_9.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_1__0_.mem_left_track_9.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_bottom_track_1.mem_out[0:7] = 8'b10000100;
	force uut.u_efpga.FPGA.sb_1__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b01111011;
	force uut.u_efpga.FPGA.sb_1__1_.mem_bottom_track_9.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_bottom_track_9.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__1_.mem_left_track_9.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_1__1_.mem_left_track_9.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_1__2_.mem_right_track_0.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__2_.mem_right_track_0.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__2_.mem_right_track_8.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_1__2_.mem_right_track_8.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_1__2_.mem_left_track_1.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__2_.mem_left_track_1.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_1__2_.mem_left_track_9.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_1__2_.mem_left_track_9.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_0.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_0.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_4.mem_out[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_9.mem_out[0:1] = 2'b10;
	force uut.u_efpga.FPGA.sb_2__0_.mem_left_track_9.mem_outb[0:1] = 2'b01;
	force uut.u_efpga.FPGA.sb_2__1_.mem_top_track_0.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_2__1_.mem_top_track_0.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_2__1_.mem_top_track_8.mem_out[0:5] = 6'b001001;
	force uut.u_efpga.FPGA.sb_2__1_.mem_top_track_8.mem_outb[0:5] = 6'b110110;
	force uut.u_efpga.FPGA.sb_2__1_.mem_bottom_track_1.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_2__1_.mem_bottom_track_1.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_2__1_.mem_bottom_track_9.mem_out[0:7] = 8'b00000001;
	force uut.u_efpga.FPGA.sb_2__1_.mem_bottom_track_9.mem_outb[0:7] = 8'b11111110;
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_7.mem_out[0:1] = 2'b01;
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_7.mem_outb[0:1] = 2'b10;
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__1_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_1.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_1.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_1.mem_out[0:5] = 6'b000001;
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_1.mem_outb[0:5] = 6'b111110;
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.sb_2__2_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_bottom_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__0_.mem_top_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__1_.mem_top_ipin_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_bottom_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_1__2_.mem_top_ipin_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_4.mem_out[0:1] = 2'b01;
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_4.mem_outb[0:1] = 2'b10;
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_bottom_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_2.mem_out[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__0_.mem_top_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_bottom_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__1_.mem_top_ipin_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_bottom_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_8.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cbx_2__2_.mem_top_ipin_8.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_left_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__1_.mem_right_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_left_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_0__2_.mem_right_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_left_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__1_.mem_right_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_left_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_1__2_.mem_right_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_left_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__1_.mem_right_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_left_ipin_7.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_0.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_0.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_1.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_1.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_2.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_2.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_3.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_3.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_4.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_4.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_5.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_5.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_6.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_6.mem_outb[0:1] = {2{1'b1}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_7.mem_out[0:1] = {2{1'b0}};
	force uut.u_efpga.FPGA.cby_2__2_.mem_right_ipin_7.mem_outb[0:1] = {2{1'b1}};
end

W25Q256JVxIQ u_spi_host_model(
.CLK  (cio_sck_o),
.CSn  (cio_csb_o),
.DIO  (cio_mosi_o),
.WPn,
.HOLDn,
.DO   (cio_miso_i)
);

always begin
#5 clk_in1 <= ~clk_in1;
end
initial begin
clk_in1 <= 0;
rst_ni <= 0;
uart_rx_i <=1;
sram_rx_i <=1;
#100 
rst_ni <= 1;
#3000us 
repeat(100) #104us  sram_rx_i <= ~sram_rx_i;

end


endmodule
