// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register slice conforming to Comportibility guide.

module prim_subreg
  import prim_subreg_pkg::*;
#(
  parameter int            DW       = 32,
  parameter sw_access_e    SwAccess = SwAccessRW,
  parameter logic [DW-1:0] RESVAL   = '0    // reset value
) (
  input clk_i,
  input rst_ni,

  // From SW: valid for RW, WO, W1C, W1S, W0C, RC
  // In case of RC, Top connects Read Pulse to we
  input          we,
  input [DW-1:0] wd,

  // From HW: valid for HRW, HWO
  input          de,
  input [DW-1:0] d,

  // output to HW and Reg Read
  output logic          qe,
  output logic [DW-1:0] q,
  output logic [DW-1:0] qs
);

  logic          wr_en;
  logic [DW-1:0] wr_data;

  prim_subreg_arb #(
    .DW       ( DW       ),
    .SwAccess ( SwAccess )
  ) wr_en_data_arb (
    .we,
    .wd,
    .de,
    .d,
    .q,
    .wr_en,
    .wr_data
  );

  always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
      qe <= 1'b0;
    end else begin
      qe <= we;
    end
  end

  logic wr_en_buf;
  prim_generic_buf #(
    .Width(1)
  ) u_wr_en_buf (
    .in_i(wr_en),
    .out_o(wr_en_buf)
  );

  always_ff @(posedge clk_i) begin
    if (!rst_ni) begin
      q <= RESVAL;
    end else if (wr_en_buf) begin
      q <= wr_data;
    end
  end

  logic [DW-1:0] q_buf;
  prim_generic_buf #(
    .Width(DW)
  ) u_q_buf (
    .in_i(q),
    .out_o(q_buf)
  );

  assign qs = q_buf;

endmodule
