`timescale 1ns / 1ps

module bitstream
#(
	parameter BITSTREAM_LENGTH = 1
)
(
	input		[$clog2(BITSTREAM_LENGTH):0]	addrRd,
	output	reg	[0:0]							dataRd
);

always @(*) begin

	case(addrRd)
       0		:	dataRd	 = 	 1'b1
;       1		:	dataRd	 = 	 1'b0
;       2		:	dataRd	 = 	 1'b0
;       3		:	dataRd	 = 	 1'b0
;       4		:	dataRd	 = 	 1'b0
;       5		:	dataRd	 = 	 1'b0
;       6		:	dataRd	 = 	 1'b0
;       7		:	dataRd	 = 	 1'b0
;       8		:	dataRd	 = 	 1'b0
;       9		:	dataRd	 = 	 1'b0
;      10		:	dataRd	 = 	 1'b0
;      11		:	dataRd	 = 	 1'b0
;      12		:	dataRd	 = 	 1'b0
;      13		:	dataRd	 = 	 1'b0
;      14		:	dataRd	 = 	 1'b0
;      15		:	dataRd	 = 	 1'b0
;      16		:	dataRd	 = 	 1'b1
;      17		:	dataRd	 = 	 1'b0
;      18		:	dataRd	 = 	 1'b0
;      19		:	dataRd	 = 	 1'b0
;      20		:	dataRd	 = 	 1'b0
;      21		:	dataRd	 = 	 1'b0
;      22		:	dataRd	 = 	 1'b0
;      23		:	dataRd	 = 	 1'b0
;      24		:	dataRd	 = 	 1'b0
;      25		:	dataRd	 = 	 1'b0
;      26		:	dataRd	 = 	 1'b0
;      27		:	dataRd	 = 	 1'b0
;      28		:	dataRd	 = 	 1'b0
;      29		:	dataRd	 = 	 1'b0
;      30		:	dataRd	 = 	 1'b0
;      31		:	dataRd	 = 	 1'b0
;      32		:	dataRd	 = 	 1'b1
;      33		:	dataRd	 = 	 1'b0
;      34		:	dataRd	 = 	 1'b0
;      35		:	dataRd	 = 	 1'b0
;      36		:	dataRd	 = 	 1'b0
;      37		:	dataRd	 = 	 1'b0
;      38		:	dataRd	 = 	 1'b0
;      39		:	dataRd	 = 	 1'b0
;      40		:	dataRd	 = 	 1'b0
;      41		:	dataRd	 = 	 1'b0
;      42		:	dataRd	 = 	 1'b0
;      43		:	dataRd	 = 	 1'b0
;      44		:	dataRd	 = 	 1'b0
;      45		:	dataRd	 = 	 1'b0
;      46		:	dataRd	 = 	 1'b0
;      47		:	dataRd	 = 	 1'b0
;      48		:	dataRd	 = 	 1'b1
;      49		:	dataRd	 = 	 1'b0
;      50		:	dataRd	 = 	 1'b0
;      51		:	dataRd	 = 	 1'b0
;      52		:	dataRd	 = 	 1'b0
;      53		:	dataRd	 = 	 1'b0
;      54		:	dataRd	 = 	 1'b0
;      55		:	dataRd	 = 	 1'b0
;      56		:	dataRd	 = 	 1'b0
;      57		:	dataRd	 = 	 1'b0
;      58		:	dataRd	 = 	 1'b0
;      59		:	dataRd	 = 	 1'b0
;      60		:	dataRd	 = 	 1'b0
;      61		:	dataRd	 = 	 1'b0
;      62		:	dataRd	 = 	 1'b0
;      63		:	dataRd	 = 	 1'b0
;      64		:	dataRd	 = 	 1'b1
;      65		:	dataRd	 = 	 1'b0
;      66		:	dataRd	 = 	 1'b0
;      67		:	dataRd	 = 	 1'b0
;      68		:	dataRd	 = 	 1'b0
;      69		:	dataRd	 = 	 1'b0
;      70		:	dataRd	 = 	 1'b0
;      71		:	dataRd	 = 	 1'b0
;      72		:	dataRd	 = 	 1'b0
;      73		:	dataRd	 = 	 1'b0
;      74		:	dataRd	 = 	 1'b0
;      75		:	dataRd	 = 	 1'b0
;      76		:	dataRd	 = 	 1'b0
;      77		:	dataRd	 = 	 1'b0
;      78		:	dataRd	 = 	 1'b0
;      79		:	dataRd	 = 	 1'b0
;      80		:	dataRd	 = 	 1'b1
;      81		:	dataRd	 = 	 1'b0
;      82		:	dataRd	 = 	 1'b0
;      83		:	dataRd	 = 	 1'b0
;      84		:	dataRd	 = 	 1'b0
;      85		:	dataRd	 = 	 1'b0
;      86		:	dataRd	 = 	 1'b0
;      87		:	dataRd	 = 	 1'b0
;      88		:	dataRd	 = 	 1'b0
;      89		:	dataRd	 = 	 1'b0
;      90		:	dataRd	 = 	 1'b0
;      91		:	dataRd	 = 	 1'b0
;      92		:	dataRd	 = 	 1'b0
;      93		:	dataRd	 = 	 1'b0
;      94		:	dataRd	 = 	 1'b0
;      95		:	dataRd	 = 	 1'b0
;      96		:	dataRd	 = 	 1'b1
;      97		:	dataRd	 = 	 1'b0
;      98		:	dataRd	 = 	 1'b0
;      99		:	dataRd	 = 	 1'b0
;     100		:	dataRd	 = 	 1'b0
;     101		:	dataRd	 = 	 1'b0
;     102		:	dataRd	 = 	 1'b0
;     103		:	dataRd	 = 	 1'b0
;     104		:	dataRd	 = 	 1'b0
;     105		:	dataRd	 = 	 1'b0
;     106		:	dataRd	 = 	 1'b0
;     107		:	dataRd	 = 	 1'b0
;     108		:	dataRd	 = 	 1'b0
;     109		:	dataRd	 = 	 1'b0
;     110		:	dataRd	 = 	 1'b0
;     111		:	dataRd	 = 	 1'b0
;     112		:	dataRd	 = 	 1'b1
;     113		:	dataRd	 = 	 1'b0
;     114		:	dataRd	 = 	 1'b0
;     115		:	dataRd	 = 	 1'b0
;     116		:	dataRd	 = 	 1'b0
;     117		:	dataRd	 = 	 1'b0
;     118		:	dataRd	 = 	 1'b0
;     119		:	dataRd	 = 	 1'b0
;     120		:	dataRd	 = 	 1'b0
;     121		:	dataRd	 = 	 1'b0
;     122		:	dataRd	 = 	 1'b0
;     123		:	dataRd	 = 	 1'b0
;     124		:	dataRd	 = 	 1'b0
;     125		:	dataRd	 = 	 1'b0
;     126		:	dataRd	 = 	 1'b0
;     127		:	dataRd	 = 	 1'b0
;     128		:	dataRd	 = 	 1'b1
;     129		:	dataRd	 = 	 1'b0
;     130		:	dataRd	 = 	 1'b0
;     131		:	dataRd	 = 	 1'b0
;     132		:	dataRd	 = 	 1'b0
;     133		:	dataRd	 = 	 1'b0
;     134		:	dataRd	 = 	 1'b0
;     135		:	dataRd	 = 	 1'b0
;     136		:	dataRd	 = 	 1'b0
;     137		:	dataRd	 = 	 1'b0
;     138		:	dataRd	 = 	 1'b0
;     139		:	dataRd	 = 	 1'b0
;     140		:	dataRd	 = 	 1'b0
;     141		:	dataRd	 = 	 1'b0
;     142		:	dataRd	 = 	 1'b0
;     143		:	dataRd	 = 	 1'b0
;     144		:	dataRd	 = 	 1'b1
;     145		:	dataRd	 = 	 1'b0
;     146		:	dataRd	 = 	 1'b0
;     147		:	dataRd	 = 	 1'b0
;     148		:	dataRd	 = 	 1'b0
;     149		:	dataRd	 = 	 1'b0
;     150		:	dataRd	 = 	 1'b0
;     151		:	dataRd	 = 	 1'b0
;     152		:	dataRd	 = 	 1'b0
;     153		:	dataRd	 = 	 1'b0
;     154		:	dataRd	 = 	 1'b0
;     155		:	dataRd	 = 	 1'b0
;     156		:	dataRd	 = 	 1'b0
;     157		:	dataRd	 = 	 1'b0
;     158		:	dataRd	 = 	 1'b0
;     159		:	dataRd	 = 	 1'b0
;     160		:	dataRd	 = 	 1'b1
;     161		:	dataRd	 = 	 1'b0
;     162		:	dataRd	 = 	 1'b0
;     163		:	dataRd	 = 	 1'b0
;     164		:	dataRd	 = 	 1'b0
;     165		:	dataRd	 = 	 1'b0
;     166		:	dataRd	 = 	 1'b0
;     167		:	dataRd	 = 	 1'b0
;     168		:	dataRd	 = 	 1'b0
;     169		:	dataRd	 = 	 1'b0
;     170		:	dataRd	 = 	 1'b0
;     171		:	dataRd	 = 	 1'b0
;     172		:	dataRd	 = 	 1'b0
;     173		:	dataRd	 = 	 1'b0
;     174		:	dataRd	 = 	 1'b0
;     175		:	dataRd	 = 	 1'b0
;     176		:	dataRd	 = 	 1'b1
;     177		:	dataRd	 = 	 1'b0
;     178		:	dataRd	 = 	 1'b0
;     179		:	dataRd	 = 	 1'b0
;     180		:	dataRd	 = 	 1'b0
;     181		:	dataRd	 = 	 1'b0
;     182		:	dataRd	 = 	 1'b0
;     183		:	dataRd	 = 	 1'b0
;     184		:	dataRd	 = 	 1'b0
;     185		:	dataRd	 = 	 1'b0
;     186		:	dataRd	 = 	 1'b0
;     187		:	dataRd	 = 	 1'b0
;     188		:	dataRd	 = 	 1'b0
;     189		:	dataRd	 = 	 1'b0
;     190		:	dataRd	 = 	 1'b0
;     191		:	dataRd	 = 	 1'b0
;     192		:	dataRd	 = 	 1'b1
;     193		:	dataRd	 = 	 1'b0
;     194		:	dataRd	 = 	 1'b0
;     195		:	dataRd	 = 	 1'b0
;     196		:	dataRd	 = 	 1'b0
;     197		:	dataRd	 = 	 1'b0
;     198		:	dataRd	 = 	 1'b0
;     199		:	dataRd	 = 	 1'b0
;     200		:	dataRd	 = 	 1'b0
;     201		:	dataRd	 = 	 1'b0
;     202		:	dataRd	 = 	 1'b0
;     203		:	dataRd	 = 	 1'b0
;     204		:	dataRd	 = 	 1'b0
;     205		:	dataRd	 = 	 1'b0
;     206		:	dataRd	 = 	 1'b0
;     207		:	dataRd	 = 	 1'b0
;     208		:	dataRd	 = 	 1'b1
;     209		:	dataRd	 = 	 1'b0
;     210		:	dataRd	 = 	 1'b0
;     211		:	dataRd	 = 	 1'b0
;     212		:	dataRd	 = 	 1'b0
;     213		:	dataRd	 = 	 1'b0
;     214		:	dataRd	 = 	 1'b0
;     215		:	dataRd	 = 	 1'b0
;     216		:	dataRd	 = 	 1'b0
;     217		:	dataRd	 = 	 1'b0
;     218		:	dataRd	 = 	 1'b0
;     219		:	dataRd	 = 	 1'b0
;     220		:	dataRd	 = 	 1'b0
;     221		:	dataRd	 = 	 1'b0
;     222		:	dataRd	 = 	 1'b0
;     223		:	dataRd	 = 	 1'b0
;     224		:	dataRd	 = 	 1'b1
;     225		:	dataRd	 = 	 1'b0
;     226		:	dataRd	 = 	 1'b0
;     227		:	dataRd	 = 	 1'b0
;     228		:	dataRd	 = 	 1'b0
;     229		:	dataRd	 = 	 1'b0
;     230		:	dataRd	 = 	 1'b0
;     231		:	dataRd	 = 	 1'b0
;     232		:	dataRd	 = 	 1'b0
;     233		:	dataRd	 = 	 1'b0
;     234		:	dataRd	 = 	 1'b0
;     235		:	dataRd	 = 	 1'b0
;     236		:	dataRd	 = 	 1'b0
;     237		:	dataRd	 = 	 1'b0
;     238		:	dataRd	 = 	 1'b0
;     239		:	dataRd	 = 	 1'b0
;     240		:	dataRd	 = 	 1'b1
;     241		:	dataRd	 = 	 1'b0
;     242		:	dataRd	 = 	 1'b0
;     243		:	dataRd	 = 	 1'b0
;     244		:	dataRd	 = 	 1'b0
;     245		:	dataRd	 = 	 1'b0
;     246		:	dataRd	 = 	 1'b0
;     247		:	dataRd	 = 	 1'b0
;     248		:	dataRd	 = 	 1'b0
;     249		:	dataRd	 = 	 1'b0
;     250		:	dataRd	 = 	 1'b0
;     251		:	dataRd	 = 	 1'b0
;     252		:	dataRd	 = 	 1'b0
;     253		:	dataRd	 = 	 1'b0
;     254		:	dataRd	 = 	 1'b0
;     255		:	dataRd	 = 	 1'b0
;     256		:	dataRd	 = 	 1'b1
;     257		:	dataRd	 = 	 1'b0
;     258		:	dataRd	 = 	 1'b0
;     259		:	dataRd	 = 	 1'b0
;     260		:	dataRd	 = 	 1'b0
;     261		:	dataRd	 = 	 1'b0
;     262		:	dataRd	 = 	 1'b0
;     263		:	dataRd	 = 	 1'b0
;     264		:	dataRd	 = 	 1'b0
;     265		:	dataRd	 = 	 1'b0
;     266		:	dataRd	 = 	 1'b0
;     267		:	dataRd	 = 	 1'b0
;     268		:	dataRd	 = 	 1'b0
;     269		:	dataRd	 = 	 1'b0
;     270		:	dataRd	 = 	 1'b0
;     271		:	dataRd	 = 	 1'b0
;     272		:	dataRd	 = 	 1'b1
;     273		:	dataRd	 = 	 1'b0
;     274		:	dataRd	 = 	 1'b0
;     275		:	dataRd	 = 	 1'b0
;     276		:	dataRd	 = 	 1'b0
;     277		:	dataRd	 = 	 1'b0
;     278		:	dataRd	 = 	 1'b0
;     279		:	dataRd	 = 	 1'b0
;     280		:	dataRd	 = 	 1'b0
;     281		:	dataRd	 = 	 1'b0
;     282		:	dataRd	 = 	 1'b0
;     283		:	dataRd	 = 	 1'b0
;     284		:	dataRd	 = 	 1'b0
;     285		:	dataRd	 = 	 1'b0
;     286		:	dataRd	 = 	 1'b0
;     287		:	dataRd	 = 	 1'b0
;     288		:	dataRd	 = 	 1'b1
;     289		:	dataRd	 = 	 1'b0
;     290		:	dataRd	 = 	 1'b0
;     291		:	dataRd	 = 	 1'b0
;     292		:	dataRd	 = 	 1'b0
;     293		:	dataRd	 = 	 1'b0
;     294		:	dataRd	 = 	 1'b0
;     295		:	dataRd	 = 	 1'b0
;     296		:	dataRd	 = 	 1'b0
;     297		:	dataRd	 = 	 1'b0
;     298		:	dataRd	 = 	 1'b0
;     299		:	dataRd	 = 	 1'b0
;     300		:	dataRd	 = 	 1'b0
;     301		:	dataRd	 = 	 1'b0
;     302		:	dataRd	 = 	 1'b0
;     303		:	dataRd	 = 	 1'b0
;     304		:	dataRd	 = 	 1'b1
;     305		:	dataRd	 = 	 1'b0
;     306		:	dataRd	 = 	 1'b0
;     307		:	dataRd	 = 	 1'b0
;     308		:	dataRd	 = 	 1'b0
;     309		:	dataRd	 = 	 1'b0
;     310		:	dataRd	 = 	 1'b0
;     311		:	dataRd	 = 	 1'b0
;     312		:	dataRd	 = 	 1'b0
;     313		:	dataRd	 = 	 1'b0
;     314		:	dataRd	 = 	 1'b0
;     315		:	dataRd	 = 	 1'b0
;     316		:	dataRd	 = 	 1'b0
;     317		:	dataRd	 = 	 1'b0
;     318		:	dataRd	 = 	 1'b0
;     319		:	dataRd	 = 	 1'b0
;     320		:	dataRd	 = 	 1'b1
;     321		:	dataRd	 = 	 1'b0
;     322		:	dataRd	 = 	 1'b0
;     323		:	dataRd	 = 	 1'b0
;     324		:	dataRd	 = 	 1'b0
;     325		:	dataRd	 = 	 1'b0
;     326		:	dataRd	 = 	 1'b0
;     327		:	dataRd	 = 	 1'b0
;     328		:	dataRd	 = 	 1'b0
;     329		:	dataRd	 = 	 1'b0
;     330		:	dataRd	 = 	 1'b0
;     331		:	dataRd	 = 	 1'b0
;     332		:	dataRd	 = 	 1'b0
;     333		:	dataRd	 = 	 1'b0
;     334		:	dataRd	 = 	 1'b0
;     335		:	dataRd	 = 	 1'b0
;     336		:	dataRd	 = 	 1'b1
;     337		:	dataRd	 = 	 1'b0
;     338		:	dataRd	 = 	 1'b0
;     339		:	dataRd	 = 	 1'b0
;     340		:	dataRd	 = 	 1'b0
;     341		:	dataRd	 = 	 1'b0
;     342		:	dataRd	 = 	 1'b0
;     343		:	dataRd	 = 	 1'b0
;     344		:	dataRd	 = 	 1'b0
;     345		:	dataRd	 = 	 1'b0
;     346		:	dataRd	 = 	 1'b0
;     347		:	dataRd	 = 	 1'b0
;     348		:	dataRd	 = 	 1'b0
;     349		:	dataRd	 = 	 1'b0
;     350		:	dataRd	 = 	 1'b0
;     351		:	dataRd	 = 	 1'b0
;     352		:	dataRd	 = 	 1'b1
;     353		:	dataRd	 = 	 1'b0
;     354		:	dataRd	 = 	 1'b0
;     355		:	dataRd	 = 	 1'b0
;     356		:	dataRd	 = 	 1'b0
;     357		:	dataRd	 = 	 1'b0
;     358		:	dataRd	 = 	 1'b0
;     359		:	dataRd	 = 	 1'b0
;     360		:	dataRd	 = 	 1'b0
;     361		:	dataRd	 = 	 1'b0
;     362		:	dataRd	 = 	 1'b0
;     363		:	dataRd	 = 	 1'b0
;     364		:	dataRd	 = 	 1'b0
;     365		:	dataRd	 = 	 1'b0
;     366		:	dataRd	 = 	 1'b0
;     367		:	dataRd	 = 	 1'b0
;     368		:	dataRd	 = 	 1'b1
;     369		:	dataRd	 = 	 1'b0
;     370		:	dataRd	 = 	 1'b0
;     371		:	dataRd	 = 	 1'b0
;     372		:	dataRd	 = 	 1'b0
;     373		:	dataRd	 = 	 1'b0
;     374		:	dataRd	 = 	 1'b0
;     375		:	dataRd	 = 	 1'b0
;     376		:	dataRd	 = 	 1'b0
;     377		:	dataRd	 = 	 1'b0
;     378		:	dataRd	 = 	 1'b0
;     379		:	dataRd	 = 	 1'b0
;     380		:	dataRd	 = 	 1'b0
;     381		:	dataRd	 = 	 1'b0
;     382		:	dataRd	 = 	 1'b0
;     383		:	dataRd	 = 	 1'b0
;     384		:	dataRd	 = 	 1'b1
;     385		:	dataRd	 = 	 1'b0
;     386		:	dataRd	 = 	 1'b0
;     387		:	dataRd	 = 	 1'b0
;     388		:	dataRd	 = 	 1'b0
;     389		:	dataRd	 = 	 1'b0
;     390		:	dataRd	 = 	 1'b0
;     391		:	dataRd	 = 	 1'b0
;     392		:	dataRd	 = 	 1'b0
;     393		:	dataRd	 = 	 1'b0
;     394		:	dataRd	 = 	 1'b0
;     395		:	dataRd	 = 	 1'b0
;     396		:	dataRd	 = 	 1'b0
;     397		:	dataRd	 = 	 1'b0
;     398		:	dataRd	 = 	 1'b0
;     399		:	dataRd	 = 	 1'b0
;     400		:	dataRd	 = 	 1'b1
;     401		:	dataRd	 = 	 1'b0
;     402		:	dataRd	 = 	 1'b0
;     403		:	dataRd	 = 	 1'b0
;     404		:	dataRd	 = 	 1'b0
;     405		:	dataRd	 = 	 1'b0
;     406		:	dataRd	 = 	 1'b0
;     407		:	dataRd	 = 	 1'b0
;     408		:	dataRd	 = 	 1'b0
;     409		:	dataRd	 = 	 1'b0
;     410		:	dataRd	 = 	 1'b0
;     411		:	dataRd	 = 	 1'b0
;     412		:	dataRd	 = 	 1'b0
;     413		:	dataRd	 = 	 1'b0
;     414		:	dataRd	 = 	 1'b0
;     415		:	dataRd	 = 	 1'b0
;     416		:	dataRd	 = 	 1'b1
;     417		:	dataRd	 = 	 1'b0
;     418		:	dataRd	 = 	 1'b0
;     419		:	dataRd	 = 	 1'b0
;     420		:	dataRd	 = 	 1'b0
;     421		:	dataRd	 = 	 1'b0
;     422		:	dataRd	 = 	 1'b0
;     423		:	dataRd	 = 	 1'b0
;     424		:	dataRd	 = 	 1'b0
;     425		:	dataRd	 = 	 1'b0
;     426		:	dataRd	 = 	 1'b0
;     427		:	dataRd	 = 	 1'b0
;     428		:	dataRd	 = 	 1'b0
;     429		:	dataRd	 = 	 1'b0
;     430		:	dataRd	 = 	 1'b0
;     431		:	dataRd	 = 	 1'b0
;     432		:	dataRd	 = 	 1'b1
;     433		:	dataRd	 = 	 1'b0
;     434		:	dataRd	 = 	 1'b0
;     435		:	dataRd	 = 	 1'b0
;     436		:	dataRd	 = 	 1'b0
;     437		:	dataRd	 = 	 1'b0
;     438		:	dataRd	 = 	 1'b0
;     439		:	dataRd	 = 	 1'b0
;     440		:	dataRd	 = 	 1'b0
;     441		:	dataRd	 = 	 1'b0
;     442		:	dataRd	 = 	 1'b0
;     443		:	dataRd	 = 	 1'b0
;     444		:	dataRd	 = 	 1'b0
;     445		:	dataRd	 = 	 1'b0
;     446		:	dataRd	 = 	 1'b0
;     447		:	dataRd	 = 	 1'b0
;     448		:	dataRd	 = 	 1'b1
;     449		:	dataRd	 = 	 1'b0
;     450		:	dataRd	 = 	 1'b0
;     451		:	dataRd	 = 	 1'b0
;     452		:	dataRd	 = 	 1'b0
;     453		:	dataRd	 = 	 1'b0
;     454		:	dataRd	 = 	 1'b0
;     455		:	dataRd	 = 	 1'b0
;     456		:	dataRd	 = 	 1'b0
;     457		:	dataRd	 = 	 1'b0
;     458		:	dataRd	 = 	 1'b0
;     459		:	dataRd	 = 	 1'b0
;     460		:	dataRd	 = 	 1'b0
;     461		:	dataRd	 = 	 1'b0
;     462		:	dataRd	 = 	 1'b0
;     463		:	dataRd	 = 	 1'b0
;     464		:	dataRd	 = 	 1'b1
;     465		:	dataRd	 = 	 1'b0
;     466		:	dataRd	 = 	 1'b0
;     467		:	dataRd	 = 	 1'b0
;     468		:	dataRd	 = 	 1'b0
;     469		:	dataRd	 = 	 1'b0
;     470		:	dataRd	 = 	 1'b0
;     471		:	dataRd	 = 	 1'b0
;     472		:	dataRd	 = 	 1'b0
;     473		:	dataRd	 = 	 1'b0
;     474		:	dataRd	 = 	 1'b0
;     475		:	dataRd	 = 	 1'b0
;     476		:	dataRd	 = 	 1'b0
;     477		:	dataRd	 = 	 1'b0
;     478		:	dataRd	 = 	 1'b0
;     479		:	dataRd	 = 	 1'b0
;     480		:	dataRd	 = 	 1'b1
;     481		:	dataRd	 = 	 1'b0
;     482		:	dataRd	 = 	 1'b0
;     483		:	dataRd	 = 	 1'b0
;     484		:	dataRd	 = 	 1'b0
;     485		:	dataRd	 = 	 1'b0
;     486		:	dataRd	 = 	 1'b0
;     487		:	dataRd	 = 	 1'b0
;     488		:	dataRd	 = 	 1'b0
;     489		:	dataRd	 = 	 1'b0
;     490		:	dataRd	 = 	 1'b0
;     491		:	dataRd	 = 	 1'b0
;     492		:	dataRd	 = 	 1'b0
;     493		:	dataRd	 = 	 1'b0
;     494		:	dataRd	 = 	 1'b0
;     495		:	dataRd	 = 	 1'b0
;     496		:	dataRd	 = 	 1'b1
;     497		:	dataRd	 = 	 1'b0
;     498		:	dataRd	 = 	 1'b0
;     499		:	dataRd	 = 	 1'b0
;     500		:	dataRd	 = 	 1'b0
;     501		:	dataRd	 = 	 1'b0
;     502		:	dataRd	 = 	 1'b0
;     503		:	dataRd	 = 	 1'b0
;     504		:	dataRd	 = 	 1'b0
;     505		:	dataRd	 = 	 1'b0
;     506		:	dataRd	 = 	 1'b0
;     507		:	dataRd	 = 	 1'b0
;     508		:	dataRd	 = 	 1'b0
;     509		:	dataRd	 = 	 1'b0
;     510		:	dataRd	 = 	 1'b0
;     511		:	dataRd	 = 	 1'b0
;     512		:	dataRd	 = 	 1'b1
;     513		:	dataRd	 = 	 1'b0
;     514		:	dataRd	 = 	 1'b0
;     515		:	dataRd	 = 	 1'b0
;     516		:	dataRd	 = 	 1'b0
;     517		:	dataRd	 = 	 1'b0
;     518		:	dataRd	 = 	 1'b0
;     519		:	dataRd	 = 	 1'b0
;     520		:	dataRd	 = 	 1'b0
;     521		:	dataRd	 = 	 1'b0
;     522		:	dataRd	 = 	 1'b0
;     523		:	dataRd	 = 	 1'b0
;     524		:	dataRd	 = 	 1'b0
;     525		:	dataRd	 = 	 1'b0
;     526		:	dataRd	 = 	 1'b0
;     527		:	dataRd	 = 	 1'b0
;     528		:	dataRd	 = 	 1'b1
;     529		:	dataRd	 = 	 1'b0
;     530		:	dataRd	 = 	 1'b0
;     531		:	dataRd	 = 	 1'b0
;     532		:	dataRd	 = 	 1'b0
;     533		:	dataRd	 = 	 1'b0
;     534		:	dataRd	 = 	 1'b0
;     535		:	dataRd	 = 	 1'b0
;     536		:	dataRd	 = 	 1'b0
;     537		:	dataRd	 = 	 1'b0
;     538		:	dataRd	 = 	 1'b0
;     539		:	dataRd	 = 	 1'b0
;     540		:	dataRd	 = 	 1'b0
;     541		:	dataRd	 = 	 1'b0
;     542		:	dataRd	 = 	 1'b0
;     543		:	dataRd	 = 	 1'b0
;     544		:	dataRd	 = 	 1'b1
;     545		:	dataRd	 = 	 1'b0
;     546		:	dataRd	 = 	 1'b0
;     547		:	dataRd	 = 	 1'b0
;     548		:	dataRd	 = 	 1'b0
;     549		:	dataRd	 = 	 1'b0
;     550		:	dataRd	 = 	 1'b0
;     551		:	dataRd	 = 	 1'b0
;     552		:	dataRd	 = 	 1'b0
;     553		:	dataRd	 = 	 1'b0
;     554		:	dataRd	 = 	 1'b0
;     555		:	dataRd	 = 	 1'b0
;     556		:	dataRd	 = 	 1'b0
;     557		:	dataRd	 = 	 1'b0
;     558		:	dataRd	 = 	 1'b0
;     559		:	dataRd	 = 	 1'b0
;     560		:	dataRd	 = 	 1'b1
;     561		:	dataRd	 = 	 1'b0
;     562		:	dataRd	 = 	 1'b0
;     563		:	dataRd	 = 	 1'b0
;     564		:	dataRd	 = 	 1'b0
;     565		:	dataRd	 = 	 1'b0
;     566		:	dataRd	 = 	 1'b0
;     567		:	dataRd	 = 	 1'b0
;     568		:	dataRd	 = 	 1'b0
;     569		:	dataRd	 = 	 1'b0
;     570		:	dataRd	 = 	 1'b0
;     571		:	dataRd	 = 	 1'b0
;     572		:	dataRd	 = 	 1'b0
;     573		:	dataRd	 = 	 1'b0
;     574		:	dataRd	 = 	 1'b0
;     575		:	dataRd	 = 	 1'b0
;     576		:	dataRd	 = 	 1'b1
;     577		:	dataRd	 = 	 1'b0
;     578		:	dataRd	 = 	 1'b0
;     579		:	dataRd	 = 	 1'b0
;     580		:	dataRd	 = 	 1'b0
;     581		:	dataRd	 = 	 1'b0
;     582		:	dataRd	 = 	 1'b0
;     583		:	dataRd	 = 	 1'b0
;     584		:	dataRd	 = 	 1'b0
;     585		:	dataRd	 = 	 1'b0
;     586		:	dataRd	 = 	 1'b0
;     587		:	dataRd	 = 	 1'b0
;     588		:	dataRd	 = 	 1'b0
;     589		:	dataRd	 = 	 1'b0
;     590		:	dataRd	 = 	 1'b0
;     591		:	dataRd	 = 	 1'b0
;     592		:	dataRd	 = 	 1'b1
;     593		:	dataRd	 = 	 1'b0
;     594		:	dataRd	 = 	 1'b0
;     595		:	dataRd	 = 	 1'b0
;     596		:	dataRd	 = 	 1'b0
;     597		:	dataRd	 = 	 1'b0
;     598		:	dataRd	 = 	 1'b0
;     599		:	dataRd	 = 	 1'b0
;     600		:	dataRd	 = 	 1'b0
;     601		:	dataRd	 = 	 1'b0
;     602		:	dataRd	 = 	 1'b0
;     603		:	dataRd	 = 	 1'b0
;     604		:	dataRd	 = 	 1'b0
;     605		:	dataRd	 = 	 1'b0
;     606		:	dataRd	 = 	 1'b0
;     607		:	dataRd	 = 	 1'b0
;     608		:	dataRd	 = 	 1'b1
;     609		:	dataRd	 = 	 1'b0
;     610		:	dataRd	 = 	 1'b0
;     611		:	dataRd	 = 	 1'b0
;     612		:	dataRd	 = 	 1'b0
;     613		:	dataRd	 = 	 1'b0
;     614		:	dataRd	 = 	 1'b0
;     615		:	dataRd	 = 	 1'b0
;     616		:	dataRd	 = 	 1'b0
;     617		:	dataRd	 = 	 1'b0
;     618		:	dataRd	 = 	 1'b0
;     619		:	dataRd	 = 	 1'b0
;     620		:	dataRd	 = 	 1'b0
;     621		:	dataRd	 = 	 1'b0
;     622		:	dataRd	 = 	 1'b0
;     623		:	dataRd	 = 	 1'b0
;     624		:	dataRd	 = 	 1'b1
;     625		:	dataRd	 = 	 1'b0
;     626		:	dataRd	 = 	 1'b0
;     627		:	dataRd	 = 	 1'b0
;     628		:	dataRd	 = 	 1'b0
;     629		:	dataRd	 = 	 1'b0
;     630		:	dataRd	 = 	 1'b0
;     631		:	dataRd	 = 	 1'b0
;     632		:	dataRd	 = 	 1'b0
;     633		:	dataRd	 = 	 1'b0
;     634		:	dataRd	 = 	 1'b0
;     635		:	dataRd	 = 	 1'b0
;     636		:	dataRd	 = 	 1'b0
;     637		:	dataRd	 = 	 1'b0
;     638		:	dataRd	 = 	 1'b0
;     639		:	dataRd	 = 	 1'b0
;     640		:	dataRd	 = 	 1'b1
;     641		:	dataRd	 = 	 1'b0
;     642		:	dataRd	 = 	 1'b0
;     643		:	dataRd	 = 	 1'b0
;     644		:	dataRd	 = 	 1'b0
;     645		:	dataRd	 = 	 1'b0
;     646		:	dataRd	 = 	 1'b0
;     647		:	dataRd	 = 	 1'b0
;     648		:	dataRd	 = 	 1'b0
;     649		:	dataRd	 = 	 1'b0
;     650		:	dataRd	 = 	 1'b0
;     651		:	dataRd	 = 	 1'b0
;     652		:	dataRd	 = 	 1'b0
;     653		:	dataRd	 = 	 1'b0
;     654		:	dataRd	 = 	 1'b0
;     655		:	dataRd	 = 	 1'b0
;     656		:	dataRd	 = 	 1'b1
;     657		:	dataRd	 = 	 1'b0
;     658		:	dataRd	 = 	 1'b0
;     659		:	dataRd	 = 	 1'b0
;     660		:	dataRd	 = 	 1'b0
;     661		:	dataRd	 = 	 1'b0
;     662		:	dataRd	 = 	 1'b0
;     663		:	dataRd	 = 	 1'b0
;     664		:	dataRd	 = 	 1'b0
;     665		:	dataRd	 = 	 1'b0
;     666		:	dataRd	 = 	 1'b0
;     667		:	dataRd	 = 	 1'b0
;     668		:	dataRd	 = 	 1'b0
;     669		:	dataRd	 = 	 1'b0
;     670		:	dataRd	 = 	 1'b0
;     671		:	dataRd	 = 	 1'b0
;     672		:	dataRd	 = 	 1'b1
;     673		:	dataRd	 = 	 1'b0
;     674		:	dataRd	 = 	 1'b0
;     675		:	dataRd	 = 	 1'b0
;     676		:	dataRd	 = 	 1'b0
;     677		:	dataRd	 = 	 1'b0
;     678		:	dataRd	 = 	 1'b0
;     679		:	dataRd	 = 	 1'b0
;     680		:	dataRd	 = 	 1'b0
;     681		:	dataRd	 = 	 1'b0
;     682		:	dataRd	 = 	 1'b0
;     683		:	dataRd	 = 	 1'b0
;     684		:	dataRd	 = 	 1'b0
;     685		:	dataRd	 = 	 1'b0
;     686		:	dataRd	 = 	 1'b0
;     687		:	dataRd	 = 	 1'b0
;     688		:	dataRd	 = 	 1'b1
;     689		:	dataRd	 = 	 1'b0
;     690		:	dataRd	 = 	 1'b0
;     691		:	dataRd	 = 	 1'b0
;     692		:	dataRd	 = 	 1'b0
;     693		:	dataRd	 = 	 1'b0
;     694		:	dataRd	 = 	 1'b0
;     695		:	dataRd	 = 	 1'b0
;     696		:	dataRd	 = 	 1'b0
;     697		:	dataRd	 = 	 1'b0
;     698		:	dataRd	 = 	 1'b0
;     699		:	dataRd	 = 	 1'b0
;     700		:	dataRd	 = 	 1'b0
;     701		:	dataRd	 = 	 1'b0
;     702		:	dataRd	 = 	 1'b0
;     703		:	dataRd	 = 	 1'b0
;     704		:	dataRd	 = 	 1'b1
;     705		:	dataRd	 = 	 1'b0
;     706		:	dataRd	 = 	 1'b0
;     707		:	dataRd	 = 	 1'b0
;     708		:	dataRd	 = 	 1'b0
;     709		:	dataRd	 = 	 1'b0
;     710		:	dataRd	 = 	 1'b0
;     711		:	dataRd	 = 	 1'b0
;     712		:	dataRd	 = 	 1'b0
;     713		:	dataRd	 = 	 1'b0
;     714		:	dataRd	 = 	 1'b0
;     715		:	dataRd	 = 	 1'b0
;     716		:	dataRd	 = 	 1'b0
;     717		:	dataRd	 = 	 1'b0
;     718		:	dataRd	 = 	 1'b0
;     719		:	dataRd	 = 	 1'b0
;     720		:	dataRd	 = 	 1'b1
;     721		:	dataRd	 = 	 1'b0
;     722		:	dataRd	 = 	 1'b0
;     723		:	dataRd	 = 	 1'b0
;     724		:	dataRd	 = 	 1'b0
;     725		:	dataRd	 = 	 1'b0
;     726		:	dataRd	 = 	 1'b0
;     727		:	dataRd	 = 	 1'b0
;     728		:	dataRd	 = 	 1'b0
;     729		:	dataRd	 = 	 1'b0
;     730		:	dataRd	 = 	 1'b0
;     731		:	dataRd	 = 	 1'b0
;     732		:	dataRd	 = 	 1'b0
;     733		:	dataRd	 = 	 1'b0
;     734		:	dataRd	 = 	 1'b0
;     735		:	dataRd	 = 	 1'b0
;     736		:	dataRd	 = 	 1'b1
;     737		:	dataRd	 = 	 1'b0
;     738		:	dataRd	 = 	 1'b0
;     739		:	dataRd	 = 	 1'b0
;     740		:	dataRd	 = 	 1'b0
;     741		:	dataRd	 = 	 1'b0
;     742		:	dataRd	 = 	 1'b0
;     743		:	dataRd	 = 	 1'b0
;     744		:	dataRd	 = 	 1'b0
;     745		:	dataRd	 = 	 1'b0
;     746		:	dataRd	 = 	 1'b0
;     747		:	dataRd	 = 	 1'b0
;     748		:	dataRd	 = 	 1'b0
;     749		:	dataRd	 = 	 1'b0
;     750		:	dataRd	 = 	 1'b0
;     751		:	dataRd	 = 	 1'b0
;     752		:	dataRd	 = 	 1'b1
;     753		:	dataRd	 = 	 1'b0
;     754		:	dataRd	 = 	 1'b0
;     755		:	dataRd	 = 	 1'b0
;     756		:	dataRd	 = 	 1'b0
;     757		:	dataRd	 = 	 1'b0
;     758		:	dataRd	 = 	 1'b0
;     759		:	dataRd	 = 	 1'b0
;     760		:	dataRd	 = 	 1'b0
;     761		:	dataRd	 = 	 1'b0
;     762		:	dataRd	 = 	 1'b0
;     763		:	dataRd	 = 	 1'b0
;     764		:	dataRd	 = 	 1'b0
;     765		:	dataRd	 = 	 1'b0
;     766		:	dataRd	 = 	 1'b0
;     767		:	dataRd	 = 	 1'b0
;     768		:	dataRd	 = 	 1'b1
;     769		:	dataRd	 = 	 1'b0
;     770		:	dataRd	 = 	 1'b0
;     771		:	dataRd	 = 	 1'b0
;     772		:	dataRd	 = 	 1'b0
;     773		:	dataRd	 = 	 1'b0
;     774		:	dataRd	 = 	 1'b0
;     775		:	dataRd	 = 	 1'b0
;     776		:	dataRd	 = 	 1'b0
;     777		:	dataRd	 = 	 1'b0
;     778		:	dataRd	 = 	 1'b0
;     779		:	dataRd	 = 	 1'b0
;     780		:	dataRd	 = 	 1'b0
;     781		:	dataRd	 = 	 1'b0
;     782		:	dataRd	 = 	 1'b0
;     783		:	dataRd	 = 	 1'b0
;     784		:	dataRd	 = 	 1'b1
;     785		:	dataRd	 = 	 1'b0
;     786		:	dataRd	 = 	 1'b0
;     787		:	dataRd	 = 	 1'b0
;     788		:	dataRd	 = 	 1'b0
;     789		:	dataRd	 = 	 1'b0
;     790		:	dataRd	 = 	 1'b0
;     791		:	dataRd	 = 	 1'b0
;     792		:	dataRd	 = 	 1'b0
;     793		:	dataRd	 = 	 1'b0
;     794		:	dataRd	 = 	 1'b0
;     795		:	dataRd	 = 	 1'b0
;     796		:	dataRd	 = 	 1'b0
;     797		:	dataRd	 = 	 1'b0
;     798		:	dataRd	 = 	 1'b0
;     799		:	dataRd	 = 	 1'b0
;     800		:	dataRd	 = 	 1'b1
;     801		:	dataRd	 = 	 1'b0
;     802		:	dataRd	 = 	 1'b0
;     803		:	dataRd	 = 	 1'b0
;     804		:	dataRd	 = 	 1'b0
;     805		:	dataRd	 = 	 1'b0
;     806		:	dataRd	 = 	 1'b0
;     807		:	dataRd	 = 	 1'b0
;     808		:	dataRd	 = 	 1'b0
;     809		:	dataRd	 = 	 1'b0
;     810		:	dataRd	 = 	 1'b0
;     811		:	dataRd	 = 	 1'b0
;     812		:	dataRd	 = 	 1'b0
;     813		:	dataRd	 = 	 1'b0
;     814		:	dataRd	 = 	 1'b0
;     815		:	dataRd	 = 	 1'b0
;     816		:	dataRd	 = 	 1'b1
;     817		:	dataRd	 = 	 1'b0
;     818		:	dataRd	 = 	 1'b0
;     819		:	dataRd	 = 	 1'b0
;     820		:	dataRd	 = 	 1'b0
;     821		:	dataRd	 = 	 1'b0
;     822		:	dataRd	 = 	 1'b0
;     823		:	dataRd	 = 	 1'b0
;     824		:	dataRd	 = 	 1'b0
;     825		:	dataRd	 = 	 1'b0
;     826		:	dataRd	 = 	 1'b0
;     827		:	dataRd	 = 	 1'b0
;     828		:	dataRd	 = 	 1'b0
;     829		:	dataRd	 = 	 1'b0
;     830		:	dataRd	 = 	 1'b0
;     831		:	dataRd	 = 	 1'b0
;     832		:	dataRd	 = 	 1'b1
;     833		:	dataRd	 = 	 1'b0
;     834		:	dataRd	 = 	 1'b0
;     835		:	dataRd	 = 	 1'b0
;     836		:	dataRd	 = 	 1'b0
;     837		:	dataRd	 = 	 1'b0
;     838		:	dataRd	 = 	 1'b0
;     839		:	dataRd	 = 	 1'b0
;     840		:	dataRd	 = 	 1'b0
;     841		:	dataRd	 = 	 1'b0
;     842		:	dataRd	 = 	 1'b0
;     843		:	dataRd	 = 	 1'b0
;     844		:	dataRd	 = 	 1'b0
;     845		:	dataRd	 = 	 1'b0
;     846		:	dataRd	 = 	 1'b0
;     847		:	dataRd	 = 	 1'b0
;     848		:	dataRd	 = 	 1'b1
;     849		:	dataRd	 = 	 1'b0
;     850		:	dataRd	 = 	 1'b0
;     851		:	dataRd	 = 	 1'b0
;     852		:	dataRd	 = 	 1'b0
;     853		:	dataRd	 = 	 1'b0
;     854		:	dataRd	 = 	 1'b0
;     855		:	dataRd	 = 	 1'b0
;     856		:	dataRd	 = 	 1'b0
;     857		:	dataRd	 = 	 1'b0
;     858		:	dataRd	 = 	 1'b0
;     859		:	dataRd	 = 	 1'b0
;     860		:	dataRd	 = 	 1'b0
;     861		:	dataRd	 = 	 1'b0
;     862		:	dataRd	 = 	 1'b0
;     863		:	dataRd	 = 	 1'b0
;     864		:	dataRd	 = 	 1'b1
;     865		:	dataRd	 = 	 1'b0
;     866		:	dataRd	 = 	 1'b0
;     867		:	dataRd	 = 	 1'b0
;     868		:	dataRd	 = 	 1'b0
;     869		:	dataRd	 = 	 1'b0
;     870		:	dataRd	 = 	 1'b0
;     871		:	dataRd	 = 	 1'b0
;     872		:	dataRd	 = 	 1'b0
;     873		:	dataRd	 = 	 1'b0
;     874		:	dataRd	 = 	 1'b0
;     875		:	dataRd	 = 	 1'b0
;     876		:	dataRd	 = 	 1'b0
;     877		:	dataRd	 = 	 1'b0
;     878		:	dataRd	 = 	 1'b0
;     879		:	dataRd	 = 	 1'b0
;     880		:	dataRd	 = 	 1'b1
;     881		:	dataRd	 = 	 1'b0
;     882		:	dataRd	 = 	 1'b0
;     883		:	dataRd	 = 	 1'b0
;     884		:	dataRd	 = 	 1'b0
;     885		:	dataRd	 = 	 1'b0
;     886		:	dataRd	 = 	 1'b0
;     887		:	dataRd	 = 	 1'b0
;     888		:	dataRd	 = 	 1'b0
;     889		:	dataRd	 = 	 1'b0
;     890		:	dataRd	 = 	 1'b0
;     891		:	dataRd	 = 	 1'b0
;     892		:	dataRd	 = 	 1'b0
;     893		:	dataRd	 = 	 1'b0
;     894		:	dataRd	 = 	 1'b0
;     895		:	dataRd	 = 	 1'b0
;     896		:	dataRd	 = 	 1'b1
;     897		:	dataRd	 = 	 1'b0
;     898		:	dataRd	 = 	 1'b0
;     899		:	dataRd	 = 	 1'b0
;     900		:	dataRd	 = 	 1'b0
;     901		:	dataRd	 = 	 1'b0
;     902		:	dataRd	 = 	 1'b0
;     903		:	dataRd	 = 	 1'b0
;     904		:	dataRd	 = 	 1'b0
;     905		:	dataRd	 = 	 1'b0
;     906		:	dataRd	 = 	 1'b0
;     907		:	dataRd	 = 	 1'b0
;     908		:	dataRd	 = 	 1'b0
;     909		:	dataRd	 = 	 1'b0
;     910		:	dataRd	 = 	 1'b0
;     911		:	dataRd	 = 	 1'b0
;     912		:	dataRd	 = 	 1'b1
;     913		:	dataRd	 = 	 1'b0
;     914		:	dataRd	 = 	 1'b0
;     915		:	dataRd	 = 	 1'b0
;     916		:	dataRd	 = 	 1'b0
;     917		:	dataRd	 = 	 1'b0
;     918		:	dataRd	 = 	 1'b0
;     919		:	dataRd	 = 	 1'b0
;     920		:	dataRd	 = 	 1'b0
;     921		:	dataRd	 = 	 1'b0
;     922		:	dataRd	 = 	 1'b0
;     923		:	dataRd	 = 	 1'b0
;     924		:	dataRd	 = 	 1'b0
;     925		:	dataRd	 = 	 1'b0
;     926		:	dataRd	 = 	 1'b0
;     927		:	dataRd	 = 	 1'b0
;     928		:	dataRd	 = 	 1'b1
;     929		:	dataRd	 = 	 1'b0
;     930		:	dataRd	 = 	 1'b0
;     931		:	dataRd	 = 	 1'b0
;     932		:	dataRd	 = 	 1'b0
;     933		:	dataRd	 = 	 1'b0
;     934		:	dataRd	 = 	 1'b0
;     935		:	dataRd	 = 	 1'b0
;     936		:	dataRd	 = 	 1'b0
;     937		:	dataRd	 = 	 1'b0
;     938		:	dataRd	 = 	 1'b0
;     939		:	dataRd	 = 	 1'b0
;     940		:	dataRd	 = 	 1'b0
;     941		:	dataRd	 = 	 1'b0
;     942		:	dataRd	 = 	 1'b0
;     943		:	dataRd	 = 	 1'b0
;     944		:	dataRd	 = 	 1'b1
;     945		:	dataRd	 = 	 1'b0
;     946		:	dataRd	 = 	 1'b0
;     947		:	dataRd	 = 	 1'b0
;     948		:	dataRd	 = 	 1'b0
;     949		:	dataRd	 = 	 1'b0
;     950		:	dataRd	 = 	 1'b0
;     951		:	dataRd	 = 	 1'b0
;     952		:	dataRd	 = 	 1'b0
;     953		:	dataRd	 = 	 1'b0
;     954		:	dataRd	 = 	 1'b0
;     955		:	dataRd	 = 	 1'b0
;     956		:	dataRd	 = 	 1'b0
;     957		:	dataRd	 = 	 1'b0
;     958		:	dataRd	 = 	 1'b0
;     959		:	dataRd	 = 	 1'b0
;     960		:	dataRd	 = 	 1'b1
;     961		:	dataRd	 = 	 1'b0
;     962		:	dataRd	 = 	 1'b0
;     963		:	dataRd	 = 	 1'b0
;     964		:	dataRd	 = 	 1'b0
;     965		:	dataRd	 = 	 1'b0
;     966		:	dataRd	 = 	 1'b0
;     967		:	dataRd	 = 	 1'b0
;     968		:	dataRd	 = 	 1'b0
;     969		:	dataRd	 = 	 1'b0
;     970		:	dataRd	 = 	 1'b0
;     971		:	dataRd	 = 	 1'b0
;     972		:	dataRd	 = 	 1'b0
;     973		:	dataRd	 = 	 1'b0
;     974		:	dataRd	 = 	 1'b0
;     975		:	dataRd	 = 	 1'b0
;     976		:	dataRd	 = 	 1'b0
;     977		:	dataRd	 = 	 1'b0
;     978		:	dataRd	 = 	 1'b0
;     979		:	dataRd	 = 	 1'b0
;     980		:	dataRd	 = 	 1'b0
;     981		:	dataRd	 = 	 1'b0
;     982		:	dataRd	 = 	 1'b0
;     983		:	dataRd	 = 	 1'b0
;     984		:	dataRd	 = 	 1'b0
;     985		:	dataRd	 = 	 1'b0
;     986		:	dataRd	 = 	 1'b0
;     987		:	dataRd	 = 	 1'b0
;     988		:	dataRd	 = 	 1'b0
;     989		:	dataRd	 = 	 1'b0
;     990		:	dataRd	 = 	 1'b0
;     991		:	dataRd	 = 	 1'b0
;     992		:	dataRd	 = 	 1'b0
;     993		:	dataRd	 = 	 1'b0
;     994		:	dataRd	 = 	 1'b0
;     995		:	dataRd	 = 	 1'b0
;     996		:	dataRd	 = 	 1'b0
;     997		:	dataRd	 = 	 1'b0
;     998		:	dataRd	 = 	 1'b0
;     999		:	dataRd	 = 	 1'b0
;    1000		:	dataRd	 = 	 1'b0
;    1001		:	dataRd	 = 	 1'b0
;    1002		:	dataRd	 = 	 1'b0
;    1003		:	dataRd	 = 	 1'b0
;    1004		:	dataRd	 = 	 1'b0
;    1005		:	dataRd	 = 	 1'b0
;    1006		:	dataRd	 = 	 1'b0
;    1007		:	dataRd	 = 	 1'b0
;    1008		:	dataRd	 = 	 1'b0
;    1009		:	dataRd	 = 	 1'b0
;    1010		:	dataRd	 = 	 1'b0
;    1011		:	dataRd	 = 	 1'b0
;    1012		:	dataRd	 = 	 1'b0
;    1013		:	dataRd	 = 	 1'b0
;    1014		:	dataRd	 = 	 1'b0
;    1015		:	dataRd	 = 	 1'b0
;    1016		:	dataRd	 = 	 1'b0
;    1017		:	dataRd	 = 	 1'b0
;    1018		:	dataRd	 = 	 1'b0
;    1019		:	dataRd	 = 	 1'b0
;    1020		:	dataRd	 = 	 1'b0
;    1021		:	dataRd	 = 	 1'b0
;    1022		:	dataRd	 = 	 1'b0
;    1023		:	dataRd	 = 	 1'b0
;    1024		:	dataRd	 = 	 1'b0
;    1025		:	dataRd	 = 	 1'b0
;    1026		:	dataRd	 = 	 1'b0
;    1027		:	dataRd	 = 	 1'b1
;    1028		:	dataRd	 = 	 1'b0
;    1029		:	dataRd	 = 	 1'b0
;    1030		:	dataRd	 = 	 1'b0
;    1031		:	dataRd	 = 	 1'b0
;    1032		:	dataRd	 = 	 1'b0
;    1033		:	dataRd	 = 	 1'b0
;    1034		:	dataRd	 = 	 1'b0
;    1035		:	dataRd	 = 	 1'b0
;    1036		:	dataRd	 = 	 1'b0
;    1037		:	dataRd	 = 	 1'b0
;    1038		:	dataRd	 = 	 1'b0
;    1039		:	dataRd	 = 	 1'b0
;    1040		:	dataRd	 = 	 1'b0
;    1041		:	dataRd	 = 	 1'b0
;    1042		:	dataRd	 = 	 1'b0
;    1043		:	dataRd	 = 	 1'b0
;    1044		:	dataRd	 = 	 1'b0
;    1045		:	dataRd	 = 	 1'b0
;    1046		:	dataRd	 = 	 1'b0
;    1047		:	dataRd	 = 	 1'b0
;    1048		:	dataRd	 = 	 1'b0
;    1049		:	dataRd	 = 	 1'b0
;    1050		:	dataRd	 = 	 1'b0
;    1051		:	dataRd	 = 	 1'b0
;    1052		:	dataRd	 = 	 1'b0
;    1053		:	dataRd	 = 	 1'b0
;    1054		:	dataRd	 = 	 1'b0
;    1055		:	dataRd	 = 	 1'b0
;    1056		:	dataRd	 = 	 1'b0
;    1057		:	dataRd	 = 	 1'b0
;    1058		:	dataRd	 = 	 1'b0
;    1059		:	dataRd	 = 	 1'b0
;    1060		:	dataRd	 = 	 1'b0
;    1061		:	dataRd	 = 	 1'b0
;    1062		:	dataRd	 = 	 1'b0
;    1063		:	dataRd	 = 	 1'b0
;    1064		:	dataRd	 = 	 1'b0
;    1065		:	dataRd	 = 	 1'b0
;    1066		:	dataRd	 = 	 1'b0
;    1067		:	dataRd	 = 	 1'b0
;    1068		:	dataRd	 = 	 1'b0
;    1069		:	dataRd	 = 	 1'b0
;    1070		:	dataRd	 = 	 1'b0
;    1071		:	dataRd	 = 	 1'b0
;    1072		:	dataRd	 = 	 1'b0
;    1073		:	dataRd	 = 	 1'b0
;    1074		:	dataRd	 = 	 1'b0
;    1075		:	dataRd	 = 	 1'b0
;    1076		:	dataRd	 = 	 1'b0
;    1077		:	dataRd	 = 	 1'b0
;    1078		:	dataRd	 = 	 1'b0
;    1079		:	dataRd	 = 	 1'b0
;    1080		:	dataRd	 = 	 1'b0
;    1081		:	dataRd	 = 	 1'b0
;    1082		:	dataRd	 = 	 1'b0
;    1083		:	dataRd	 = 	 1'b0
;    1084		:	dataRd	 = 	 1'b0
;    1085		:	dataRd	 = 	 1'b0
;    1086		:	dataRd	 = 	 1'b0
;    1087		:	dataRd	 = 	 1'b0
;    1088		:	dataRd	 = 	 1'b0
;    1089		:	dataRd	 = 	 1'b0
;    1090		:	dataRd	 = 	 1'b0
;    1091		:	dataRd	 = 	 1'b0
;    1092		:	dataRd	 = 	 1'b0
;    1093		:	dataRd	 = 	 1'b0
;    1094		:	dataRd	 = 	 1'b1
;    1095		:	dataRd	 = 	 1'b0
;    1096		:	dataRd	 = 	 1'b0
;    1097		:	dataRd	 = 	 1'b0
;    1098		:	dataRd	 = 	 1'b0
;    1099		:	dataRd	 = 	 1'b0
;    1100		:	dataRd	 = 	 1'b0
;    1101		:	dataRd	 = 	 1'b0
;    1102		:	dataRd	 = 	 1'b0
;    1103		:	dataRd	 = 	 1'b0
;    1104		:	dataRd	 = 	 1'b0
;    1105		:	dataRd	 = 	 1'b0
;    1106		:	dataRd	 = 	 1'b0
;    1107		:	dataRd	 = 	 1'b0
;    1108		:	dataRd	 = 	 1'b0
;    1109		:	dataRd	 = 	 1'b0
;    1110		:	dataRd	 = 	 1'b0
;    1111		:	dataRd	 = 	 1'b0
;    1112		:	dataRd	 = 	 1'b0
;    1113		:	dataRd	 = 	 1'b0
;    1114		:	dataRd	 = 	 1'b0
;    1115		:	dataRd	 = 	 1'b0
;    1116		:	dataRd	 = 	 1'b0
;    1117		:	dataRd	 = 	 1'b0
;    1118		:	dataRd	 = 	 1'b0
;    1119		:	dataRd	 = 	 1'b0
;    1120		:	dataRd	 = 	 1'b0
;    1121		:	dataRd	 = 	 1'b0
;    1122		:	dataRd	 = 	 1'b0
;    1123		:	dataRd	 = 	 1'b0
;    1124		:	dataRd	 = 	 1'b0
;    1125		:	dataRd	 = 	 1'b0
;    1126		:	dataRd	 = 	 1'b0
;    1127		:	dataRd	 = 	 1'b0
;    1128		:	dataRd	 = 	 1'b0
;    1129		:	dataRd	 = 	 1'b0
;    1130		:	dataRd	 = 	 1'b0
;    1131		:	dataRd	 = 	 1'b0
;    1132		:	dataRd	 = 	 1'b0
;    1133		:	dataRd	 = 	 1'b0
;    1134		:	dataRd	 = 	 1'b0
;    1135		:	dataRd	 = 	 1'b0
;    1136		:	dataRd	 = 	 1'b0
;    1137		:	dataRd	 = 	 1'b0
;    1138		:	dataRd	 = 	 1'b0
;    1139		:	dataRd	 = 	 1'b0
;    1140		:	dataRd	 = 	 1'b0
;    1141		:	dataRd	 = 	 1'b0
;    1142		:	dataRd	 = 	 1'b0
;    1143		:	dataRd	 = 	 1'b0
;    1144		:	dataRd	 = 	 1'b0
;    1145		:	dataRd	 = 	 1'b0
;    1146		:	dataRd	 = 	 1'b0
;    1147		:	dataRd	 = 	 1'b0
;    1148		:	dataRd	 = 	 1'b0
;    1149		:	dataRd	 = 	 1'b0
;    1150		:	dataRd	 = 	 1'b0
;    1151		:	dataRd	 = 	 1'b0
;    1152		:	dataRd	 = 	 1'b0
;    1153		:	dataRd	 = 	 1'b0
;    1154		:	dataRd	 = 	 1'b0
;    1155		:	dataRd	 = 	 1'b0
;    1156		:	dataRd	 = 	 1'b0
;    1157		:	dataRd	 = 	 1'b0
;    1158		:	dataRd	 = 	 1'b0
;    1159		:	dataRd	 = 	 1'b0
;    1160		:	dataRd	 = 	 1'b0
;    1161		:	dataRd	 = 	 1'b1
;    1162		:	dataRd	 = 	 1'b0
;    1163		:	dataRd	 = 	 1'b0
;    1164		:	dataRd	 = 	 1'b0
;    1165		:	dataRd	 = 	 1'b0
;    1166		:	dataRd	 = 	 1'b0
;    1167		:	dataRd	 = 	 1'b0
;    1168		:	dataRd	 = 	 1'b0
;    1169		:	dataRd	 = 	 1'b0
;    1170		:	dataRd	 = 	 1'b0
;    1171		:	dataRd	 = 	 1'b0
;    1172		:	dataRd	 = 	 1'b0
;    1173		:	dataRd	 = 	 1'b0
;    1174		:	dataRd	 = 	 1'b0
;    1175		:	dataRd	 = 	 1'b0
;    1176		:	dataRd	 = 	 1'b0
;    1177		:	dataRd	 = 	 1'b0
;    1178		:	dataRd	 = 	 1'b0
;    1179		:	dataRd	 = 	 1'b0
;    1180		:	dataRd	 = 	 1'b0
;    1181		:	dataRd	 = 	 1'b0
;    1182		:	dataRd	 = 	 1'b0
;    1183		:	dataRd	 = 	 1'b0
;    1184		:	dataRd	 = 	 1'b0
;    1185		:	dataRd	 = 	 1'b0
;    1186		:	dataRd	 = 	 1'b0
;    1187		:	dataRd	 = 	 1'b0
;    1188		:	dataRd	 = 	 1'b0
;    1189		:	dataRd	 = 	 1'b0
;    1190		:	dataRd	 = 	 1'b0
;    1191		:	dataRd	 = 	 1'b0
;    1192		:	dataRd	 = 	 1'b0
;    1193		:	dataRd	 = 	 1'b0
;    1194		:	dataRd	 = 	 1'b0
;    1195		:	dataRd	 = 	 1'b0
;    1196		:	dataRd	 = 	 1'b0
;    1197		:	dataRd	 = 	 1'b0
;    1198		:	dataRd	 = 	 1'b0
;    1199		:	dataRd	 = 	 1'b0
;    1200		:	dataRd	 = 	 1'b0
;    1201		:	dataRd	 = 	 1'b0
;    1202		:	dataRd	 = 	 1'b0
;    1203		:	dataRd	 = 	 1'b0
;    1204		:	dataRd	 = 	 1'b0
;    1205		:	dataRd	 = 	 1'b0
;    1206		:	dataRd	 = 	 1'b0
;    1207		:	dataRd	 = 	 1'b0
;    1208		:	dataRd	 = 	 1'b0
;    1209		:	dataRd	 = 	 1'b0
;    1210		:	dataRd	 = 	 1'b0
;    1211		:	dataRd	 = 	 1'b0
;    1212		:	dataRd	 = 	 1'b0
;    1213		:	dataRd	 = 	 1'b0
;    1214		:	dataRd	 = 	 1'b0
;    1215		:	dataRd	 = 	 1'b0
;    1216		:	dataRd	 = 	 1'b0
;    1217		:	dataRd	 = 	 1'b0
;    1218		:	dataRd	 = 	 1'b0
;    1219		:	dataRd	 = 	 1'b0
;    1220		:	dataRd	 = 	 1'b0
;    1221		:	dataRd	 = 	 1'b0
;    1222		:	dataRd	 = 	 1'b0
;    1223		:	dataRd	 = 	 1'b0
;    1224		:	dataRd	 = 	 1'b0
;    1225		:	dataRd	 = 	 1'b0
;    1226		:	dataRd	 = 	 1'b0
;    1227		:	dataRd	 = 	 1'b0
;    1228		:	dataRd	 = 	 1'b1
;    1229		:	dataRd	 = 	 1'b0
;    1230		:	dataRd	 = 	 1'b0
;    1231		:	dataRd	 = 	 1'b0
;    1232		:	dataRd	 = 	 1'b0
;    1233		:	dataRd	 = 	 1'b0
;    1234		:	dataRd	 = 	 1'b0
;    1235		:	dataRd	 = 	 1'b0
;    1236		:	dataRd	 = 	 1'b0
;    1237		:	dataRd	 = 	 1'b0
;    1238		:	dataRd	 = 	 1'b0
;    1239		:	dataRd	 = 	 1'b0
;    1240		:	dataRd	 = 	 1'b0
;    1241		:	dataRd	 = 	 1'b0
;    1242		:	dataRd	 = 	 1'b0
;    1243		:	dataRd	 = 	 1'b0
;    1244		:	dataRd	 = 	 1'b0
;    1245		:	dataRd	 = 	 1'b0
;    1246		:	dataRd	 = 	 1'b0
;    1247		:	dataRd	 = 	 1'b0
;    1248		:	dataRd	 = 	 1'b0
;    1249		:	dataRd	 = 	 1'b0
;    1250		:	dataRd	 = 	 1'b0
;    1251		:	dataRd	 = 	 1'b0
;    1252		:	dataRd	 = 	 1'b0
;    1253		:	dataRd	 = 	 1'b0
;    1254		:	dataRd	 = 	 1'b0
;    1255		:	dataRd	 = 	 1'b0
;    1256		:	dataRd	 = 	 1'b0
;    1257		:	dataRd	 = 	 1'b0
;    1258		:	dataRd	 = 	 1'b0
;    1259		:	dataRd	 = 	 1'b0
;    1260		:	dataRd	 = 	 1'b0
;    1261		:	dataRd	 = 	 1'b0
;    1262		:	dataRd	 = 	 1'b0
;    1263		:	dataRd	 = 	 1'b0
;    1264		:	dataRd	 = 	 1'b0
;    1265		:	dataRd	 = 	 1'b0
;    1266		:	dataRd	 = 	 1'b0
;    1267		:	dataRd	 = 	 1'b0
;    1268		:	dataRd	 = 	 1'b0
;    1269		:	dataRd	 = 	 1'b0
;    1270		:	dataRd	 = 	 1'b0
;    1271		:	dataRd	 = 	 1'b0
;    1272		:	dataRd	 = 	 1'b0
;    1273		:	dataRd	 = 	 1'b0
;    1274		:	dataRd	 = 	 1'b0
;    1275		:	dataRd	 = 	 1'b0
;    1276		:	dataRd	 = 	 1'b0
;    1277		:	dataRd	 = 	 1'b0
;    1278		:	dataRd	 = 	 1'b0
;    1279		:	dataRd	 = 	 1'b0
;    1280		:	dataRd	 = 	 1'b0
;    1281		:	dataRd	 = 	 1'b0
;    1282		:	dataRd	 = 	 1'b0
;    1283		:	dataRd	 = 	 1'b0
;    1284		:	dataRd	 = 	 1'b0
;    1285		:	dataRd	 = 	 1'b0
;    1286		:	dataRd	 = 	 1'b0
;    1287		:	dataRd	 = 	 1'b0
;    1288		:	dataRd	 = 	 1'b0
;    1289		:	dataRd	 = 	 1'b0
;    1290		:	dataRd	 = 	 1'b0
;    1291		:	dataRd	 = 	 1'b0
;    1292		:	dataRd	 = 	 1'b0
;    1293		:	dataRd	 = 	 1'b0
;    1294		:	dataRd	 = 	 1'b0
;    1295		:	dataRd	 = 	 1'b1
;    1296		:	dataRd	 = 	 1'b0
;    1297		:	dataRd	 = 	 1'b0
;    1298		:	dataRd	 = 	 1'b0
;    1299		:	dataRd	 = 	 1'b0
;    1300		:	dataRd	 = 	 1'b0
;    1301		:	dataRd	 = 	 1'b0
;    1302		:	dataRd	 = 	 1'b0
;    1303		:	dataRd	 = 	 1'b0
;    1304		:	dataRd	 = 	 1'b0
;    1305		:	dataRd	 = 	 1'b0
;    1306		:	dataRd	 = 	 1'b0
;    1307		:	dataRd	 = 	 1'b0
;    1308		:	dataRd	 = 	 1'b0
;    1309		:	dataRd	 = 	 1'b0
;    1310		:	dataRd	 = 	 1'b0
;    1311		:	dataRd	 = 	 1'b0
;    1312		:	dataRd	 = 	 1'b0
;    1313		:	dataRd	 = 	 1'b0
;    1314		:	dataRd	 = 	 1'b0
;    1315		:	dataRd	 = 	 1'b0
;    1316		:	dataRd	 = 	 1'b0
;    1317		:	dataRd	 = 	 1'b0
;    1318		:	dataRd	 = 	 1'b0
;    1319		:	dataRd	 = 	 1'b0
;    1320		:	dataRd	 = 	 1'b0
;    1321		:	dataRd	 = 	 1'b0
;    1322		:	dataRd	 = 	 1'b0
;    1323		:	dataRd	 = 	 1'b0
;    1324		:	dataRd	 = 	 1'b0
;    1325		:	dataRd	 = 	 1'b0
;    1326		:	dataRd	 = 	 1'b0
;    1327		:	dataRd	 = 	 1'b0
;    1328		:	dataRd	 = 	 1'b0
;    1329		:	dataRd	 = 	 1'b0
;    1330		:	dataRd	 = 	 1'b0
;    1331		:	dataRd	 = 	 1'b0
;    1332		:	dataRd	 = 	 1'b0
;    1333		:	dataRd	 = 	 1'b0
;    1334		:	dataRd	 = 	 1'b0
;    1335		:	dataRd	 = 	 1'b0
;    1336		:	dataRd	 = 	 1'b0
;    1337		:	dataRd	 = 	 1'b0
;    1338		:	dataRd	 = 	 1'b0
;    1339		:	dataRd	 = 	 1'b0
;    1340		:	dataRd	 = 	 1'b0
;    1341		:	dataRd	 = 	 1'b0
;    1342		:	dataRd	 = 	 1'b0
;    1343		:	dataRd	 = 	 1'b0
;    1344		:	dataRd	 = 	 1'b0
;    1345		:	dataRd	 = 	 1'b0
;    1346		:	dataRd	 = 	 1'b0
;    1347		:	dataRd	 = 	 1'b0
;    1348		:	dataRd	 = 	 1'b0
;    1349		:	dataRd	 = 	 1'b0
;    1350		:	dataRd	 = 	 1'b0
;    1351		:	dataRd	 = 	 1'b0
;    1352		:	dataRd	 = 	 1'b0
;    1353		:	dataRd	 = 	 1'b0
;    1354		:	dataRd	 = 	 1'b0
;    1355		:	dataRd	 = 	 1'b0
;    1356		:	dataRd	 = 	 1'b0
;    1357		:	dataRd	 = 	 1'b0
;    1358		:	dataRd	 = 	 1'b0
;    1359		:	dataRd	 = 	 1'b0
;    1360		:	dataRd	 = 	 1'b0
;    1361		:	dataRd	 = 	 1'b0
;    1362		:	dataRd	 = 	 1'b1
;    1363		:	dataRd	 = 	 1'b0
;    1364		:	dataRd	 = 	 1'b0
;    1365		:	dataRd	 = 	 1'b0
;    1366		:	dataRd	 = 	 1'b0
;    1367		:	dataRd	 = 	 1'b0
;    1368		:	dataRd	 = 	 1'b0
;    1369		:	dataRd	 = 	 1'b0
;    1370		:	dataRd	 = 	 1'b0
;    1371		:	dataRd	 = 	 1'b0
;    1372		:	dataRd	 = 	 1'b0
;    1373		:	dataRd	 = 	 1'b0
;    1374		:	dataRd	 = 	 1'b0
;    1375		:	dataRd	 = 	 1'b0
;    1376		:	dataRd	 = 	 1'b0
;    1377		:	dataRd	 = 	 1'b0
;    1378		:	dataRd	 = 	 1'b0
;    1379		:	dataRd	 = 	 1'b0
;    1380		:	dataRd	 = 	 1'b0
;    1381		:	dataRd	 = 	 1'b0
;    1382		:	dataRd	 = 	 1'b0
;    1383		:	dataRd	 = 	 1'b0
;    1384		:	dataRd	 = 	 1'b0
;    1385		:	dataRd	 = 	 1'b0
;    1386		:	dataRd	 = 	 1'b0
;    1387		:	dataRd	 = 	 1'b0
;    1388		:	dataRd	 = 	 1'b0
;    1389		:	dataRd	 = 	 1'b0
;    1390		:	dataRd	 = 	 1'b0
;    1391		:	dataRd	 = 	 1'b0
;    1392		:	dataRd	 = 	 1'b0
;    1393		:	dataRd	 = 	 1'b0
;    1394		:	dataRd	 = 	 1'b0
;    1395		:	dataRd	 = 	 1'b0
;    1396		:	dataRd	 = 	 1'b0
;    1397		:	dataRd	 = 	 1'b0
;    1398		:	dataRd	 = 	 1'b0
;    1399		:	dataRd	 = 	 1'b0
;    1400		:	dataRd	 = 	 1'b0
;    1401		:	dataRd	 = 	 1'b0
;    1402		:	dataRd	 = 	 1'b0
;    1403		:	dataRd	 = 	 1'b0
;    1404		:	dataRd	 = 	 1'b0
;    1405		:	dataRd	 = 	 1'b0
;    1406		:	dataRd	 = 	 1'b0
;    1407		:	dataRd	 = 	 1'b0
;    1408		:	dataRd	 = 	 1'b0
;    1409		:	dataRd	 = 	 1'b0
;    1410		:	dataRd	 = 	 1'b0
;    1411		:	dataRd	 = 	 1'b0
;    1412		:	dataRd	 = 	 1'b0
;    1413		:	dataRd	 = 	 1'b0
;    1414		:	dataRd	 = 	 1'b0
;    1415		:	dataRd	 = 	 1'b0
;    1416		:	dataRd	 = 	 1'b0
;    1417		:	dataRd	 = 	 1'b0
;    1418		:	dataRd	 = 	 1'b0
;    1419		:	dataRd	 = 	 1'b0
;    1420		:	dataRd	 = 	 1'b0
;    1421		:	dataRd	 = 	 1'b0
;    1422		:	dataRd	 = 	 1'b0
;    1423		:	dataRd	 = 	 1'b0
;    1424		:	dataRd	 = 	 1'b0
;    1425		:	dataRd	 = 	 1'b0
;    1426		:	dataRd	 = 	 1'b0
;    1427		:	dataRd	 = 	 1'b0
;    1428		:	dataRd	 = 	 1'b0
;    1429		:	dataRd	 = 	 1'b1
;    1430		:	dataRd	 = 	 1'b0
;    1431		:	dataRd	 = 	 1'b0
;    1432		:	dataRd	 = 	 1'b0
;    1433		:	dataRd	 = 	 1'b0
;    1434		:	dataRd	 = 	 1'b0
;    1435		:	dataRd	 = 	 1'b0
;    1436		:	dataRd	 = 	 1'b0
;    1437		:	dataRd	 = 	 1'b0
;    1438		:	dataRd	 = 	 1'b0
;    1439		:	dataRd	 = 	 1'b0
;    1440		:	dataRd	 = 	 1'b0
;    1441		:	dataRd	 = 	 1'b0
;    1442		:	dataRd	 = 	 1'b0
;    1443		:	dataRd	 = 	 1'b0
;    1444		:	dataRd	 = 	 1'b0
;    1445		:	dataRd	 = 	 1'b0
;    1446		:	dataRd	 = 	 1'b0
;    1447		:	dataRd	 = 	 1'b0
;    1448		:	dataRd	 = 	 1'b0
;    1449		:	dataRd	 = 	 1'b0
;    1450		:	dataRd	 = 	 1'b0
;    1451		:	dataRd	 = 	 1'b0
;    1452		:	dataRd	 = 	 1'b0
;    1453		:	dataRd	 = 	 1'b0
;    1454		:	dataRd	 = 	 1'b0
;    1455		:	dataRd	 = 	 1'b0
;    1456		:	dataRd	 = 	 1'b0
;    1457		:	dataRd	 = 	 1'b0
;    1458		:	dataRd	 = 	 1'b0
;    1459		:	dataRd	 = 	 1'b0
;    1460		:	dataRd	 = 	 1'b0
;    1461		:	dataRd	 = 	 1'b0
;    1462		:	dataRd	 = 	 1'b0
;    1463		:	dataRd	 = 	 1'b0
;    1464		:	dataRd	 = 	 1'b0
;    1465		:	dataRd	 = 	 1'b0
;    1466		:	dataRd	 = 	 1'b0
;    1467		:	dataRd	 = 	 1'b0
;    1468		:	dataRd	 = 	 1'b0
;    1469		:	dataRd	 = 	 1'b0
;    1470		:	dataRd	 = 	 1'b0
;    1471		:	dataRd	 = 	 1'b0
;    1472		:	dataRd	 = 	 1'b0
;    1473		:	dataRd	 = 	 1'b0
;    1474		:	dataRd	 = 	 1'b0
;    1475		:	dataRd	 = 	 1'b0
;    1476		:	dataRd	 = 	 1'b0
;    1477		:	dataRd	 = 	 1'b0
;    1478		:	dataRd	 = 	 1'b0
;    1479		:	dataRd	 = 	 1'b0
;    1480		:	dataRd	 = 	 1'b0
;    1481		:	dataRd	 = 	 1'b0
;    1482		:	dataRd	 = 	 1'b0
;    1483		:	dataRd	 = 	 1'b0
;    1484		:	dataRd	 = 	 1'b0
;    1485		:	dataRd	 = 	 1'b0
;    1486		:	dataRd	 = 	 1'b0
;    1487		:	dataRd	 = 	 1'b0
;    1488		:	dataRd	 = 	 1'b0
;    1489		:	dataRd	 = 	 1'b0
;    1490		:	dataRd	 = 	 1'b0
;    1491		:	dataRd	 = 	 1'b0
;    1492		:	dataRd	 = 	 1'b0
;    1493		:	dataRd	 = 	 1'b0
;    1494		:	dataRd	 = 	 1'b0
;    1495		:	dataRd	 = 	 1'b0
;    1496		:	dataRd	 = 	 1'b1
;    1497		:	dataRd	 = 	 1'b0
;    1498		:	dataRd	 = 	 1'b0
;    1499		:	dataRd	 = 	 1'b0
;    1500		:	dataRd	 = 	 1'b0
;    1501		:	dataRd	 = 	 1'b0
;    1502		:	dataRd	 = 	 1'b0
;    1503		:	dataRd	 = 	 1'b0
;    1504		:	dataRd	 = 	 1'b0
;    1505		:	dataRd	 = 	 1'b0
;    1506		:	dataRd	 = 	 1'b0
;    1507		:	dataRd	 = 	 1'b0
;    1508		:	dataRd	 = 	 1'b0
;    1509		:	dataRd	 = 	 1'b0
;    1510		:	dataRd	 = 	 1'b0
;    1511		:	dataRd	 = 	 1'b0
;    1512		:	dataRd	 = 	 1'b0
;    1513		:	dataRd	 = 	 1'b0
;    1514		:	dataRd	 = 	 1'b0
;    1515		:	dataRd	 = 	 1'b0
;    1516		:	dataRd	 = 	 1'b0
;    1517		:	dataRd	 = 	 1'b0
;    1518		:	dataRd	 = 	 1'b0
;    1519		:	dataRd	 = 	 1'b0
;    1520		:	dataRd	 = 	 1'b0
;    1521		:	dataRd	 = 	 1'b0
;    1522		:	dataRd	 = 	 1'b0
;    1523		:	dataRd	 = 	 1'b0
;    1524		:	dataRd	 = 	 1'b0
;    1525		:	dataRd	 = 	 1'b0
;    1526		:	dataRd	 = 	 1'b0
;    1527		:	dataRd	 = 	 1'b0
;    1528		:	dataRd	 = 	 1'b0
;    1529		:	dataRd	 = 	 1'b0
;    1530		:	dataRd	 = 	 1'b0
;    1531		:	dataRd	 = 	 1'b0
;    1532		:	dataRd	 = 	 1'b0
;    1533		:	dataRd	 = 	 1'b0
;    1534		:	dataRd	 = 	 1'b0
;    1535		:	dataRd	 = 	 1'b0
;    1536		:	dataRd	 = 	 1'b0
;    1537		:	dataRd	 = 	 1'b0
;    1538		:	dataRd	 = 	 1'b0
;    1539		:	dataRd	 = 	 1'b0
;    1540		:	dataRd	 = 	 1'b0
;    1541		:	dataRd	 = 	 1'b0
;    1542		:	dataRd	 = 	 1'b0
;    1543		:	dataRd	 = 	 1'b0
;    1544		:	dataRd	 = 	 1'b0
;    1545		:	dataRd	 = 	 1'b0
;    1546		:	dataRd	 = 	 1'b0
;    1547		:	dataRd	 = 	 1'b0
;    1548		:	dataRd	 = 	 1'b0
;    1549		:	dataRd	 = 	 1'b0
;    1550		:	dataRd	 = 	 1'b0
;    1551		:	dataRd	 = 	 1'b0
;    1552		:	dataRd	 = 	 1'b0
;    1553		:	dataRd	 = 	 1'b0
;    1554		:	dataRd	 = 	 1'b0
;    1555		:	dataRd	 = 	 1'b0
;    1556		:	dataRd	 = 	 1'b0
;    1557		:	dataRd	 = 	 1'b0
;    1558		:	dataRd	 = 	 1'b0
;    1559		:	dataRd	 = 	 1'b0
;    1560		:	dataRd	 = 	 1'b0
;    1561		:	dataRd	 = 	 1'b0
;    1562		:	dataRd	 = 	 1'b0
;    1563		:	dataRd	 = 	 1'b1
;    1564		:	dataRd	 = 	 1'b0
;    1565		:	dataRd	 = 	 1'b0
;    1566		:	dataRd	 = 	 1'b0
;    1567		:	dataRd	 = 	 1'b0
;    1568		:	dataRd	 = 	 1'b0
;    1569		:	dataRd	 = 	 1'b0
;    1570		:	dataRd	 = 	 1'b0
;    1571		:	dataRd	 = 	 1'b0
;    1572		:	dataRd	 = 	 1'b0
;    1573		:	dataRd	 = 	 1'b0
;    1574		:	dataRd	 = 	 1'b0
;    1575		:	dataRd	 = 	 1'b0
;    1576		:	dataRd	 = 	 1'b0
;    1577		:	dataRd	 = 	 1'b0
;    1578		:	dataRd	 = 	 1'b0
;    1579		:	dataRd	 = 	 1'b0
;    1580		:	dataRd	 = 	 1'b0
;    1581		:	dataRd	 = 	 1'b0
;    1582		:	dataRd	 = 	 1'b0
;    1583		:	dataRd	 = 	 1'b0
;    1584		:	dataRd	 = 	 1'b0
;    1585		:	dataRd	 = 	 1'b0
;    1586		:	dataRd	 = 	 1'b0
;    1587		:	dataRd	 = 	 1'b0
;    1588		:	dataRd	 = 	 1'b0
;    1589		:	dataRd	 = 	 1'b0
;    1590		:	dataRd	 = 	 1'b0
;    1591		:	dataRd	 = 	 1'b0
;    1592		:	dataRd	 = 	 1'b0
;    1593		:	dataRd	 = 	 1'b0
;    1594		:	dataRd	 = 	 1'b0
;    1595		:	dataRd	 = 	 1'b0
;    1596		:	dataRd	 = 	 1'b0
;    1597		:	dataRd	 = 	 1'b0
;    1598		:	dataRd	 = 	 1'b0
;    1599		:	dataRd	 = 	 1'b0
;    1600		:	dataRd	 = 	 1'b0
;    1601		:	dataRd	 = 	 1'b0
;    1602		:	dataRd	 = 	 1'b0
;    1603		:	dataRd	 = 	 1'b0
;    1604		:	dataRd	 = 	 1'b0
;    1605		:	dataRd	 = 	 1'b0
;    1606		:	dataRd	 = 	 1'b0
;    1607		:	dataRd	 = 	 1'b0
;    1608		:	dataRd	 = 	 1'b0
;    1609		:	dataRd	 = 	 1'b0
;    1610		:	dataRd	 = 	 1'b0
;    1611		:	dataRd	 = 	 1'b0
;    1612		:	dataRd	 = 	 1'b0
;    1613		:	dataRd	 = 	 1'b0
;    1614		:	dataRd	 = 	 1'b0
;    1615		:	dataRd	 = 	 1'b0
;    1616		:	dataRd	 = 	 1'b0
;    1617		:	dataRd	 = 	 1'b0
;    1618		:	dataRd	 = 	 1'b0
;    1619		:	dataRd	 = 	 1'b0
;    1620		:	dataRd	 = 	 1'b0
;    1621		:	dataRd	 = 	 1'b0
;    1622		:	dataRd	 = 	 1'b0
;    1623		:	dataRd	 = 	 1'b0
;    1624		:	dataRd	 = 	 1'b0
;    1625		:	dataRd	 = 	 1'b0
;    1626		:	dataRd	 = 	 1'b0
;    1627		:	dataRd	 = 	 1'b0
;    1628		:	dataRd	 = 	 1'b0
;    1629		:	dataRd	 = 	 1'b0
;    1630		:	dataRd	 = 	 1'b0
;    1631		:	dataRd	 = 	 1'b0
;    1632		:	dataRd	 = 	 1'b0
;    1633		:	dataRd	 = 	 1'b0
;    1634		:	dataRd	 = 	 1'b0
;    1635		:	dataRd	 = 	 1'b0
;    1636		:	dataRd	 = 	 1'b0
;    1637		:	dataRd	 = 	 1'b0
;    1638		:	dataRd	 = 	 1'b0
;    1639		:	dataRd	 = 	 1'b0
;    1640		:	dataRd	 = 	 1'b0
;    1641		:	dataRd	 = 	 1'b0
;    1642		:	dataRd	 = 	 1'b0
;    1643		:	dataRd	 = 	 1'b0
;    1644		:	dataRd	 = 	 1'b0
;    1645		:	dataRd	 = 	 1'b0
;    1646		:	dataRd	 = 	 1'b0
;    1647		:	dataRd	 = 	 1'b0
;    1648		:	dataRd	 = 	 1'b0
;    1649		:	dataRd	 = 	 1'b0
;    1650		:	dataRd	 = 	 1'b0
;    1651		:	dataRd	 = 	 1'b0
;    1652		:	dataRd	 = 	 1'b0
;    1653		:	dataRd	 = 	 1'b0
;    1654		:	dataRd	 = 	 1'b0
;    1655		:	dataRd	 = 	 1'b0
;    1656		:	dataRd	 = 	 1'b0
;    1657		:	dataRd	 = 	 1'b0
;    1658		:	dataRd	 = 	 1'b0
;    1659		:	dataRd	 = 	 1'b0
;    1660		:	dataRd	 = 	 1'b0
;    1661		:	dataRd	 = 	 1'b0
;    1662		:	dataRd	 = 	 1'b0
;    1663		:	dataRd	 = 	 1'b0
;    1664		:	dataRd	 = 	 1'b0
;    1665		:	dataRd	 = 	 1'b0
;    1666		:	dataRd	 = 	 1'b0
;    1667		:	dataRd	 = 	 1'b0
;    1668		:	dataRd	 = 	 1'b0
;    1669		:	dataRd	 = 	 1'b0
;    1670		:	dataRd	 = 	 1'b0
;    1671		:	dataRd	 = 	 1'b0
;    1672		:	dataRd	 = 	 1'b0
;    1673		:	dataRd	 = 	 1'b0
;    1674		:	dataRd	 = 	 1'b0
;    1675		:	dataRd	 = 	 1'b0
;    1676		:	dataRd	 = 	 1'b0
;    1677		:	dataRd	 = 	 1'b0
;    1678		:	dataRd	 = 	 1'b0
;    1679		:	dataRd	 = 	 1'b0
;    1680		:	dataRd	 = 	 1'b0
;    1681		:	dataRd	 = 	 1'b0
;    1682		:	dataRd	 = 	 1'b0
;    1683		:	dataRd	 = 	 1'b0
;    1684		:	dataRd	 = 	 1'b0
;    1685		:	dataRd	 = 	 1'b0
;    1686		:	dataRd	 = 	 1'b0
;    1687		:	dataRd	 = 	 1'b0
;    1688		:	dataRd	 = 	 1'b0
;    1689		:	dataRd	 = 	 1'b0
;    1690		:	dataRd	 = 	 1'b0
;    1691		:	dataRd	 = 	 1'b0
;    1692		:	dataRd	 = 	 1'b1
;    1693		:	dataRd	 = 	 1'b0
;    1694		:	dataRd	 = 	 1'b0
;    1695		:	dataRd	 = 	 1'b1
;    1696		:	dataRd	 = 	 1'b0
;    1697		:	dataRd	 = 	 1'b0
;    1698		:	dataRd	 = 	 1'b1
;    1699		:	dataRd	 = 	 1'b0
;    1700		:	dataRd	 = 	 1'b0
;    1701		:	dataRd	 = 	 1'b0
;    1702		:	dataRd	 = 	 1'b0
;    1703		:	dataRd	 = 	 1'b0
;    1704		:	dataRd	 = 	 1'b0
;    1705		:	dataRd	 = 	 1'b0
;    1706		:	dataRd	 = 	 1'b1
;    1707		:	dataRd	 = 	 1'b0
;    1708		:	dataRd	 = 	 1'b0
;    1709		:	dataRd	 = 	 1'b1
;    1710		:	dataRd	 = 	 1'b0
;    1711		:	dataRd	 = 	 1'b0
;    1712		:	dataRd	 = 	 1'b0
;    1713		:	dataRd	 = 	 1'b0
;    1714		:	dataRd	 = 	 1'b1
;    1715		:	dataRd	 = 	 1'b0
;    1716		:	dataRd	 = 	 1'b0
;    1717		:	dataRd	 = 	 1'b0
;    1718		:	dataRd	 = 	 1'b0
;    1719		:	dataRd	 = 	 1'b1
;    1720		:	dataRd	 = 	 1'b1
;    1721		:	dataRd	 = 	 1'b0
;    1722		:	dataRd	 = 	 1'b0
;    1723		:	dataRd	 = 	 1'b1
;    1724		:	dataRd	 = 	 1'b0
;    1725		:	dataRd	 = 	 1'b0
;    1726		:	dataRd	 = 	 1'b1
;    1727		:	dataRd	 = 	 1'b0
;    1728		:	dataRd	 = 	 1'b0
;    1729		:	dataRd	 = 	 1'b0
;    1730		:	dataRd	 = 	 1'b0
;    1731		:	dataRd	 = 	 1'b0
;    1732		:	dataRd	 = 	 1'b0
;    1733		:	dataRd	 = 	 1'b0
;    1734		:	dataRd	 = 	 1'b1
;    1735		:	dataRd	 = 	 1'b0
;    1736		:	dataRd	 = 	 1'b0
;    1737		:	dataRd	 = 	 1'b1
;    1738		:	dataRd	 = 	 1'b0
;    1739		:	dataRd	 = 	 1'b0
;    1740		:	dataRd	 = 	 1'b1
;    1741		:	dataRd	 = 	 1'b0
;    1742		:	dataRd	 = 	 1'b0
;    1743		:	dataRd	 = 	 1'b0
;    1744		:	dataRd	 = 	 1'b0
;    1745		:	dataRd	 = 	 1'b0
;    1746		:	dataRd	 = 	 1'b0
;    1747		:	dataRd	 = 	 1'b0
;    1748		:	dataRd	 = 	 1'b1
;    1749		:	dataRd	 = 	 1'b0
;    1750		:	dataRd	 = 	 1'b0
;    1751		:	dataRd	 = 	 1'b0
;    1752		:	dataRd	 = 	 1'b0
;    1753		:	dataRd	 = 	 1'b0
;    1754		:	dataRd	 = 	 1'b0
;    1755		:	dataRd	 = 	 1'b0
;    1756		:	dataRd	 = 	 1'b0
;    1757		:	dataRd	 = 	 1'b0
;    1758		:	dataRd	 = 	 1'b0
;    1759		:	dataRd	 = 	 1'b0
;    1760		:	dataRd	 = 	 1'b0
;    1761		:	dataRd	 = 	 1'b0
;    1762		:	dataRd	 = 	 1'b0
;    1763		:	dataRd	 = 	 1'b0
;    1764		:	dataRd	 = 	 1'b1
;    1765		:	dataRd	 = 	 1'b0
;    1766		:	dataRd	 = 	 1'b0
;    1767		:	dataRd	 = 	 1'b0
;    1768		:	dataRd	 = 	 1'b0
;    1769		:	dataRd	 = 	 1'b0
;    1770		:	dataRd	 = 	 1'b0
;    1771		:	dataRd	 = 	 1'b0
;    1772		:	dataRd	 = 	 1'b0
;    1773		:	dataRd	 = 	 1'b0
;    1774		:	dataRd	 = 	 1'b0
;    1775		:	dataRd	 = 	 1'b0
;    1776		:	dataRd	 = 	 1'b0
;    1777		:	dataRd	 = 	 1'b0
;    1778		:	dataRd	 = 	 1'b0
;    1779		:	dataRd	 = 	 1'b0
;    1780		:	dataRd	 = 	 1'b1
;    1781		:	dataRd	 = 	 1'b0
;    1782		:	dataRd	 = 	 1'b0
;    1783		:	dataRd	 = 	 1'b0
;    1784		:	dataRd	 = 	 1'b0
;    1785		:	dataRd	 = 	 1'b0
;    1786		:	dataRd	 = 	 1'b0
;    1787		:	dataRd	 = 	 1'b0
;    1788		:	dataRd	 = 	 1'b0
;    1789		:	dataRd	 = 	 1'b0
;    1790		:	dataRd	 = 	 1'b0
;    1791		:	dataRd	 = 	 1'b0
;    1792		:	dataRd	 = 	 1'b0
;    1793		:	dataRd	 = 	 1'b0
;    1794		:	dataRd	 = 	 1'b0
;    1795		:	dataRd	 = 	 1'b0
;    1796		:	dataRd	 = 	 1'b1
;    1797		:	dataRd	 = 	 1'b0
;    1798		:	dataRd	 = 	 1'b0
;    1799		:	dataRd	 = 	 1'b0
;    1800		:	dataRd	 = 	 1'b0
;    1801		:	dataRd	 = 	 1'b0
;    1802		:	dataRd	 = 	 1'b0
;    1803		:	dataRd	 = 	 1'b0
;    1804		:	dataRd	 = 	 1'b0
;    1805		:	dataRd	 = 	 1'b0
;    1806		:	dataRd	 = 	 1'b0
;    1807		:	dataRd	 = 	 1'b0
;    1808		:	dataRd	 = 	 1'b0
;    1809		:	dataRd	 = 	 1'b0
;    1810		:	dataRd	 = 	 1'b0
;    1811		:	dataRd	 = 	 1'b0
;    1812		:	dataRd	 = 	 1'b1
;    1813		:	dataRd	 = 	 1'b0
;    1814		:	dataRd	 = 	 1'b0
;    1815		:	dataRd	 = 	 1'b0
;    1816		:	dataRd	 = 	 1'b0
;    1817		:	dataRd	 = 	 1'b0
;    1818		:	dataRd	 = 	 1'b0
;    1819		:	dataRd	 = 	 1'b0
;    1820		:	dataRd	 = 	 1'b0
;    1821		:	dataRd	 = 	 1'b0
;    1822		:	dataRd	 = 	 1'b0
;    1823		:	dataRd	 = 	 1'b0
;    1824		:	dataRd	 = 	 1'b0
;    1825		:	dataRd	 = 	 1'b0
;    1826		:	dataRd	 = 	 1'b0
;    1827		:	dataRd	 = 	 1'b0
;    1828		:	dataRd	 = 	 1'b1
;    1829		:	dataRd	 = 	 1'b0
;    1830		:	dataRd	 = 	 1'b0
;    1831		:	dataRd	 = 	 1'b0
;    1832		:	dataRd	 = 	 1'b0
;    1833		:	dataRd	 = 	 1'b0
;    1834		:	dataRd	 = 	 1'b0
;    1835		:	dataRd	 = 	 1'b0
;    1836		:	dataRd	 = 	 1'b0
;    1837		:	dataRd	 = 	 1'b0
;    1838		:	dataRd	 = 	 1'b0
;    1839		:	dataRd	 = 	 1'b0
;    1840		:	dataRd	 = 	 1'b0
;    1841		:	dataRd	 = 	 1'b0
;    1842		:	dataRd	 = 	 1'b0
;    1843		:	dataRd	 = 	 1'b0
;    1844		:	dataRd	 = 	 1'b1
;    1845		:	dataRd	 = 	 1'b0
;    1846		:	dataRd	 = 	 1'b0
;    1847		:	dataRd	 = 	 1'b0
;    1848		:	dataRd	 = 	 1'b0
;    1849		:	dataRd	 = 	 1'b0
;    1850		:	dataRd	 = 	 1'b0
;    1851		:	dataRd	 = 	 1'b0
;    1852		:	dataRd	 = 	 1'b0
;    1853		:	dataRd	 = 	 1'b0
;    1854		:	dataRd	 = 	 1'b0
;    1855		:	dataRd	 = 	 1'b0
;    1856		:	dataRd	 = 	 1'b0
;    1857		:	dataRd	 = 	 1'b0
;    1858		:	dataRd	 = 	 1'b0
;    1859		:	dataRd	 = 	 1'b0
;    1860		:	dataRd	 = 	 1'b1
;    1861		:	dataRd	 = 	 1'b0
;    1862		:	dataRd	 = 	 1'b0
;    1863		:	dataRd	 = 	 1'b0
;    1864		:	dataRd	 = 	 1'b0
;    1865		:	dataRd	 = 	 1'b0
;    1866		:	dataRd	 = 	 1'b0
;    1867		:	dataRd	 = 	 1'b0
;    1868		:	dataRd	 = 	 1'b0
;    1869		:	dataRd	 = 	 1'b0
;    1870		:	dataRd	 = 	 1'b0
;    1871		:	dataRd	 = 	 1'b0
;    1872		:	dataRd	 = 	 1'b0
;    1873		:	dataRd	 = 	 1'b0
;    1874		:	dataRd	 = 	 1'b0
;    1875		:	dataRd	 = 	 1'b0
;    1876		:	dataRd	 = 	 1'b1
;    1877		:	dataRd	 = 	 1'b0
;    1878		:	dataRd	 = 	 1'b0
;    1879		:	dataRd	 = 	 1'b0
;    1880		:	dataRd	 = 	 1'b0
;    1881		:	dataRd	 = 	 1'b0
;    1882		:	dataRd	 = 	 1'b0
;    1883		:	dataRd	 = 	 1'b0
;    1884		:	dataRd	 = 	 1'b0
;    1885		:	dataRd	 = 	 1'b0
;    1886		:	dataRd	 = 	 1'b0
;    1887		:	dataRd	 = 	 1'b0
;    1888		:	dataRd	 = 	 1'b0
;    1889		:	dataRd	 = 	 1'b0
;    1890		:	dataRd	 = 	 1'b0
;    1891		:	dataRd	 = 	 1'b0
;    1892		:	dataRd	 = 	 1'b1
;    1893		:	dataRd	 = 	 1'b0
;    1894		:	dataRd	 = 	 1'b0
;    1895		:	dataRd	 = 	 1'b0
;    1896		:	dataRd	 = 	 1'b0
;    1897		:	dataRd	 = 	 1'b0
;    1898		:	dataRd	 = 	 1'b0
;    1899		:	dataRd	 = 	 1'b0
;    1900		:	dataRd	 = 	 1'b0
;    1901		:	dataRd	 = 	 1'b0
;    1902		:	dataRd	 = 	 1'b0
;    1903		:	dataRd	 = 	 1'b0
;    1904		:	dataRd	 = 	 1'b0
;    1905		:	dataRd	 = 	 1'b0
;    1906		:	dataRd	 = 	 1'b0
;    1907		:	dataRd	 = 	 1'b0
;    1908		:	dataRd	 = 	 1'b1
;    1909		:	dataRd	 = 	 1'b0
;    1910		:	dataRd	 = 	 1'b0
;    1911		:	dataRd	 = 	 1'b0
;    1912		:	dataRd	 = 	 1'b0
;    1913		:	dataRd	 = 	 1'b0
;    1914		:	dataRd	 = 	 1'b0
;    1915		:	dataRd	 = 	 1'b0
;    1916		:	dataRd	 = 	 1'b0
;    1917		:	dataRd	 = 	 1'b0
;    1918		:	dataRd	 = 	 1'b0
;    1919		:	dataRd	 = 	 1'b0
;    1920		:	dataRd	 = 	 1'b0
;    1921		:	dataRd	 = 	 1'b0
;    1922		:	dataRd	 = 	 1'b0
;    1923		:	dataRd	 = 	 1'b0
;    1924		:	dataRd	 = 	 1'b1
;    1925		:	dataRd	 = 	 1'b0
;    1926		:	dataRd	 = 	 1'b0
;    1927		:	dataRd	 = 	 1'b0
;    1928		:	dataRd	 = 	 1'b0
;    1929		:	dataRd	 = 	 1'b0
;    1930		:	dataRd	 = 	 1'b0
;    1931		:	dataRd	 = 	 1'b0
;    1932		:	dataRd	 = 	 1'b0
;    1933		:	dataRd	 = 	 1'b0
;    1934		:	dataRd	 = 	 1'b0
;    1935		:	dataRd	 = 	 1'b0
;    1936		:	dataRd	 = 	 1'b0
;    1937		:	dataRd	 = 	 1'b0
;    1938		:	dataRd	 = 	 1'b0
;    1939		:	dataRd	 = 	 1'b0
;    1940		:	dataRd	 = 	 1'b1
;    1941		:	dataRd	 = 	 1'b0
;    1942		:	dataRd	 = 	 1'b0
;    1943		:	dataRd	 = 	 1'b0
;    1944		:	dataRd	 = 	 1'b0
;    1945		:	dataRd	 = 	 1'b0
;    1946		:	dataRd	 = 	 1'b0
;    1947		:	dataRd	 = 	 1'b0
;    1948		:	dataRd	 = 	 1'b0
;    1949		:	dataRd	 = 	 1'b0
;    1950		:	dataRd	 = 	 1'b0
;    1951		:	dataRd	 = 	 1'b0
;    1952		:	dataRd	 = 	 1'b0
;    1953		:	dataRd	 = 	 1'b0
;    1954		:	dataRd	 = 	 1'b0
;    1955		:	dataRd	 = 	 1'b0
;    1956		:	dataRd	 = 	 1'b1
;    1957		:	dataRd	 = 	 1'b0
;    1958		:	dataRd	 = 	 1'b0
;    1959		:	dataRd	 = 	 1'b0
;    1960		:	dataRd	 = 	 1'b0
;    1961		:	dataRd	 = 	 1'b0
;    1962		:	dataRd	 = 	 1'b0
;    1963		:	dataRd	 = 	 1'b0
;    1964		:	dataRd	 = 	 1'b0
;    1965		:	dataRd	 = 	 1'b0
;    1966		:	dataRd	 = 	 1'b0
;    1967		:	dataRd	 = 	 1'b0
;    1968		:	dataRd	 = 	 1'b0
;    1969		:	dataRd	 = 	 1'b0
;    1970		:	dataRd	 = 	 1'b0
;    1971		:	dataRd	 = 	 1'b0
;    1972		:	dataRd	 = 	 1'b1
;    1973		:	dataRd	 = 	 1'b0
;    1974		:	dataRd	 = 	 1'b0
;    1975		:	dataRd	 = 	 1'b0
;    1976		:	dataRd	 = 	 1'b0
;    1977		:	dataRd	 = 	 1'b0
;    1978		:	dataRd	 = 	 1'b0
;    1979		:	dataRd	 = 	 1'b0
;    1980		:	dataRd	 = 	 1'b0
;    1981		:	dataRd	 = 	 1'b0
;    1982		:	dataRd	 = 	 1'b0
;    1983		:	dataRd	 = 	 1'b0
;    1984		:	dataRd	 = 	 1'b0
;    1985		:	dataRd	 = 	 1'b0
;    1986		:	dataRd	 = 	 1'b0
;    1987		:	dataRd	 = 	 1'b0
;    1988		:	dataRd	 = 	 1'b1
;    1989		:	dataRd	 = 	 1'b0
;    1990		:	dataRd	 = 	 1'b0
;    1991		:	dataRd	 = 	 1'b0
;    1992		:	dataRd	 = 	 1'b0
;    1993		:	dataRd	 = 	 1'b0
;    1994		:	dataRd	 = 	 1'b0
;    1995		:	dataRd	 = 	 1'b0
;    1996		:	dataRd	 = 	 1'b0
;    1997		:	dataRd	 = 	 1'b0
;    1998		:	dataRd	 = 	 1'b0
;    1999		:	dataRd	 = 	 1'b0
;    2000		:	dataRd	 = 	 1'b0
;    2001		:	dataRd	 = 	 1'b0
;    2002		:	dataRd	 = 	 1'b0
;    2003		:	dataRd	 = 	 1'b0
;    2004		:	dataRd	 = 	 1'b1
;    2005		:	dataRd	 = 	 1'b0
;    2006		:	dataRd	 = 	 1'b0
;    2007		:	dataRd	 = 	 1'b0
;    2008		:	dataRd	 = 	 1'b0
;    2009		:	dataRd	 = 	 1'b0
;    2010		:	dataRd	 = 	 1'b0
;    2011		:	dataRd	 = 	 1'b0
;    2012		:	dataRd	 = 	 1'b0
;    2013		:	dataRd	 = 	 1'b0
;    2014		:	dataRd	 = 	 1'b0
;    2015		:	dataRd	 = 	 1'b0
;    2016		:	dataRd	 = 	 1'b0
;    2017		:	dataRd	 = 	 1'b0
;    2018		:	dataRd	 = 	 1'b0
;    2019		:	dataRd	 = 	 1'b0
;    2020		:	dataRd	 = 	 1'b1
;    2021		:	dataRd	 = 	 1'b0
;    2022		:	dataRd	 = 	 1'b0
;    2023		:	dataRd	 = 	 1'b0
;    2024		:	dataRd	 = 	 1'b0
;    2025		:	dataRd	 = 	 1'b0
;    2026		:	dataRd	 = 	 1'b0
;    2027		:	dataRd	 = 	 1'b0
;    2028		:	dataRd	 = 	 1'b0
;    2029		:	dataRd	 = 	 1'b0
;    2030		:	dataRd	 = 	 1'b0
;    2031		:	dataRd	 = 	 1'b0
;    2032		:	dataRd	 = 	 1'b0
;    2033		:	dataRd	 = 	 1'b0
;    2034		:	dataRd	 = 	 1'b0
;    2035		:	dataRd	 = 	 1'b0
;    2036		:	dataRd	 = 	 1'b1
;    2037		:	dataRd	 = 	 1'b0
;    2038		:	dataRd	 = 	 1'b0
;    2039		:	dataRd	 = 	 1'b0
;    2040		:	dataRd	 = 	 1'b0
;    2041		:	dataRd	 = 	 1'b0
;    2042		:	dataRd	 = 	 1'b0
;    2043		:	dataRd	 = 	 1'b0
;    2044		:	dataRd	 = 	 1'b0
;    2045		:	dataRd	 = 	 1'b0
;    2046		:	dataRd	 = 	 1'b0
;    2047		:	dataRd	 = 	 1'b0
;    2048		:	dataRd	 = 	 1'b0
;    2049		:	dataRd	 = 	 1'b0
;    2050		:	dataRd	 = 	 1'b0
;    2051		:	dataRd	 = 	 1'b0
;    2052		:	dataRd	 = 	 1'b1
;    2053		:	dataRd	 = 	 1'b0
;    2054		:	dataRd	 = 	 1'b0
;    2055		:	dataRd	 = 	 1'b0
;    2056		:	dataRd	 = 	 1'b0
;    2057		:	dataRd	 = 	 1'b0
;    2058		:	dataRd	 = 	 1'b0
;    2059		:	dataRd	 = 	 1'b0
;    2060		:	dataRd	 = 	 1'b0
;    2061		:	dataRd	 = 	 1'b0
;    2062		:	dataRd	 = 	 1'b0
;    2063		:	dataRd	 = 	 1'b0
;    2064		:	dataRd	 = 	 1'b0
;    2065		:	dataRd	 = 	 1'b0
;    2066		:	dataRd	 = 	 1'b0
;    2067		:	dataRd	 = 	 1'b0
;    2068		:	dataRd	 = 	 1'b1
;    2069		:	dataRd	 = 	 1'b0
;    2070		:	dataRd	 = 	 1'b0
;    2071		:	dataRd	 = 	 1'b0
;    2072		:	dataRd	 = 	 1'b0
;    2073		:	dataRd	 = 	 1'b0
;    2074		:	dataRd	 = 	 1'b0
;    2075		:	dataRd	 = 	 1'b0
;    2076		:	dataRd	 = 	 1'b0
;    2077		:	dataRd	 = 	 1'b0
;    2078		:	dataRd	 = 	 1'b0
;    2079		:	dataRd	 = 	 1'b0
;    2080		:	dataRd	 = 	 1'b0
;    2081		:	dataRd	 = 	 1'b0
;    2082		:	dataRd	 = 	 1'b0
;    2083		:	dataRd	 = 	 1'b0
;    2084		:	dataRd	 = 	 1'b1
;    2085		:	dataRd	 = 	 1'b0
;    2086		:	dataRd	 = 	 1'b0
;    2087		:	dataRd	 = 	 1'b0
;    2088		:	dataRd	 = 	 1'b0
;    2089		:	dataRd	 = 	 1'b0
;    2090		:	dataRd	 = 	 1'b0
;    2091		:	dataRd	 = 	 1'b0
;    2092		:	dataRd	 = 	 1'b0
;    2093		:	dataRd	 = 	 1'b0
;    2094		:	dataRd	 = 	 1'b0
;    2095		:	dataRd	 = 	 1'b0
;    2096		:	dataRd	 = 	 1'b0
;    2097		:	dataRd	 = 	 1'b0
;    2098		:	dataRd	 = 	 1'b0
;    2099		:	dataRd	 = 	 1'b0
;    2100		:	dataRd	 = 	 1'b1
;    2101		:	dataRd	 = 	 1'b0
;    2102		:	dataRd	 = 	 1'b0
;    2103		:	dataRd	 = 	 1'b0
;    2104		:	dataRd	 = 	 1'b0
;    2105		:	dataRd	 = 	 1'b0
;    2106		:	dataRd	 = 	 1'b0
;    2107		:	dataRd	 = 	 1'b0
;    2108		:	dataRd	 = 	 1'b0
;    2109		:	dataRd	 = 	 1'b0
;    2110		:	dataRd	 = 	 1'b0
;    2111		:	dataRd	 = 	 1'b0
;    2112		:	dataRd	 = 	 1'b0
;    2113		:	dataRd	 = 	 1'b0
;    2114		:	dataRd	 = 	 1'b0
;    2115		:	dataRd	 = 	 1'b0
;    2116		:	dataRd	 = 	 1'b1
;    2117		:	dataRd	 = 	 1'b0
;    2118		:	dataRd	 = 	 1'b0
;    2119		:	dataRd	 = 	 1'b0
;    2120		:	dataRd	 = 	 1'b0
;    2121		:	dataRd	 = 	 1'b0
;    2122		:	dataRd	 = 	 1'b0
;    2123		:	dataRd	 = 	 1'b0
;    2124		:	dataRd	 = 	 1'b0
;    2125		:	dataRd	 = 	 1'b0
;    2126		:	dataRd	 = 	 1'b0
;    2127		:	dataRd	 = 	 1'b0
;    2128		:	dataRd	 = 	 1'b0
;    2129		:	dataRd	 = 	 1'b0
;    2130		:	dataRd	 = 	 1'b0
;    2131		:	dataRd	 = 	 1'b0
;    2132		:	dataRd	 = 	 1'b1
;    2133		:	dataRd	 = 	 1'b0
;    2134		:	dataRd	 = 	 1'b0
;    2135		:	dataRd	 = 	 1'b0
;    2136		:	dataRd	 = 	 1'b0
;    2137		:	dataRd	 = 	 1'b0
;    2138		:	dataRd	 = 	 1'b0
;    2139		:	dataRd	 = 	 1'b0
;    2140		:	dataRd	 = 	 1'b0
;    2141		:	dataRd	 = 	 1'b0
;    2142		:	dataRd	 = 	 1'b0
;    2143		:	dataRd	 = 	 1'b0
;    2144		:	dataRd	 = 	 1'b0
;    2145		:	dataRd	 = 	 1'b0
;    2146		:	dataRd	 = 	 1'b0
;    2147		:	dataRd	 = 	 1'b0
;    2148		:	dataRd	 = 	 1'b1
;    2149		:	dataRd	 = 	 1'b0
;    2150		:	dataRd	 = 	 1'b0
;    2151		:	dataRd	 = 	 1'b0
;    2152		:	dataRd	 = 	 1'b0
;    2153		:	dataRd	 = 	 1'b0
;    2154		:	dataRd	 = 	 1'b0
;    2155		:	dataRd	 = 	 1'b0
;    2156		:	dataRd	 = 	 1'b0
;    2157		:	dataRd	 = 	 1'b0
;    2158		:	dataRd	 = 	 1'b0
;    2159		:	dataRd	 = 	 1'b0
;    2160		:	dataRd	 = 	 1'b0
;    2161		:	dataRd	 = 	 1'b0
;    2162		:	dataRd	 = 	 1'b0
;    2163		:	dataRd	 = 	 1'b0
;    2164		:	dataRd	 = 	 1'b1
;    2165		:	dataRd	 = 	 1'b0
;    2166		:	dataRd	 = 	 1'b0
;    2167		:	dataRd	 = 	 1'b0
;    2168		:	dataRd	 = 	 1'b0
;    2169		:	dataRd	 = 	 1'b0
;    2170		:	dataRd	 = 	 1'b0
;    2171		:	dataRd	 = 	 1'b0
;    2172		:	dataRd	 = 	 1'b0
;    2173		:	dataRd	 = 	 1'b0
;    2174		:	dataRd	 = 	 1'b0
;    2175		:	dataRd	 = 	 1'b0
;    2176		:	dataRd	 = 	 1'b0
;    2177		:	dataRd	 = 	 1'b0
;    2178		:	dataRd	 = 	 1'b0
;    2179		:	dataRd	 = 	 1'b0
;    2180		:	dataRd	 = 	 1'b1
;    2181		:	dataRd	 = 	 1'b0
;    2182		:	dataRd	 = 	 1'b0
;    2183		:	dataRd	 = 	 1'b0
;    2184		:	dataRd	 = 	 1'b0
;    2185		:	dataRd	 = 	 1'b0
;    2186		:	dataRd	 = 	 1'b0
;    2187		:	dataRd	 = 	 1'b0
;    2188		:	dataRd	 = 	 1'b0
;    2189		:	dataRd	 = 	 1'b0
;    2190		:	dataRd	 = 	 1'b0
;    2191		:	dataRd	 = 	 1'b0
;    2192		:	dataRd	 = 	 1'b0
;    2193		:	dataRd	 = 	 1'b0
;    2194		:	dataRd	 = 	 1'b0
;    2195		:	dataRd	 = 	 1'b0
;    2196		:	dataRd	 = 	 1'b1
;    2197		:	dataRd	 = 	 1'b0
;    2198		:	dataRd	 = 	 1'b0
;    2199		:	dataRd	 = 	 1'b0
;    2200		:	dataRd	 = 	 1'b0
;    2201		:	dataRd	 = 	 1'b0
;    2202		:	dataRd	 = 	 1'b0
;    2203		:	dataRd	 = 	 1'b0
;    2204		:	dataRd	 = 	 1'b0
;    2205		:	dataRd	 = 	 1'b0
;    2206		:	dataRd	 = 	 1'b0
;    2207		:	dataRd	 = 	 1'b0
;    2208		:	dataRd	 = 	 1'b0
;    2209		:	dataRd	 = 	 1'b0
;    2210		:	dataRd	 = 	 1'b0
;    2211		:	dataRd	 = 	 1'b0
;    2212		:	dataRd	 = 	 1'b1
;    2213		:	dataRd	 = 	 1'b0
;    2214		:	dataRd	 = 	 1'b0
;    2215		:	dataRd	 = 	 1'b0
;    2216		:	dataRd	 = 	 1'b0
;    2217		:	dataRd	 = 	 1'b0
;    2218		:	dataRd	 = 	 1'b0
;    2219		:	dataRd	 = 	 1'b0
;    2220		:	dataRd	 = 	 1'b0
;    2221		:	dataRd	 = 	 1'b0
;    2222		:	dataRd	 = 	 1'b0
;    2223		:	dataRd	 = 	 1'b0
;    2224		:	dataRd	 = 	 1'b0
;    2225		:	dataRd	 = 	 1'b0
;    2226		:	dataRd	 = 	 1'b0
;    2227		:	dataRd	 = 	 1'b0
;    2228		:	dataRd	 = 	 1'b1
;    2229		:	dataRd	 = 	 1'b0
;    2230		:	dataRd	 = 	 1'b0
;    2231		:	dataRd	 = 	 1'b0
;    2232		:	dataRd	 = 	 1'b0
;    2233		:	dataRd	 = 	 1'b0
;    2234		:	dataRd	 = 	 1'b0
;    2235		:	dataRd	 = 	 1'b0
;    2236		:	dataRd	 = 	 1'b0
;    2237		:	dataRd	 = 	 1'b0
;    2238		:	dataRd	 = 	 1'b0
;    2239		:	dataRd	 = 	 1'b0
;    2240		:	dataRd	 = 	 1'b0
;    2241		:	dataRd	 = 	 1'b0
;    2242		:	dataRd	 = 	 1'b0
;    2243		:	dataRd	 = 	 1'b0
;    2244		:	dataRd	 = 	 1'b1
;    2245		:	dataRd	 = 	 1'b0
;    2246		:	dataRd	 = 	 1'b0
;    2247		:	dataRd	 = 	 1'b0
;    2248		:	dataRd	 = 	 1'b0
;    2249		:	dataRd	 = 	 1'b0
;    2250		:	dataRd	 = 	 1'b0
;    2251		:	dataRd	 = 	 1'b0
;    2252		:	dataRd	 = 	 1'b0
;    2253		:	dataRd	 = 	 1'b0
;    2254		:	dataRd	 = 	 1'b0
;    2255		:	dataRd	 = 	 1'b0
;    2256		:	dataRd	 = 	 1'b0
;    2257		:	dataRd	 = 	 1'b0
;    2258		:	dataRd	 = 	 1'b0
;    2259		:	dataRd	 = 	 1'b0
;    2260		:	dataRd	 = 	 1'b1
;    2261		:	dataRd	 = 	 1'b0
;    2262		:	dataRd	 = 	 1'b0
;    2263		:	dataRd	 = 	 1'b0
;    2264		:	dataRd	 = 	 1'b0
;    2265		:	dataRd	 = 	 1'b0
;    2266		:	dataRd	 = 	 1'b0
;    2267		:	dataRd	 = 	 1'b0
;    2268		:	dataRd	 = 	 1'b0
;    2269		:	dataRd	 = 	 1'b0
;    2270		:	dataRd	 = 	 1'b0
;    2271		:	dataRd	 = 	 1'b0
;    2272		:	dataRd	 = 	 1'b0
;    2273		:	dataRd	 = 	 1'b0
;    2274		:	dataRd	 = 	 1'b0
;    2275		:	dataRd	 = 	 1'b0
;    2276		:	dataRd	 = 	 1'b1
;    2277		:	dataRd	 = 	 1'b0
;    2278		:	dataRd	 = 	 1'b0
;    2279		:	dataRd	 = 	 1'b0
;    2280		:	dataRd	 = 	 1'b0
;    2281		:	dataRd	 = 	 1'b0
;    2282		:	dataRd	 = 	 1'b0
;    2283		:	dataRd	 = 	 1'b0
;    2284		:	dataRd	 = 	 1'b0
;    2285		:	dataRd	 = 	 1'b0
;    2286		:	dataRd	 = 	 1'b0
;    2287		:	dataRd	 = 	 1'b0
;    2288		:	dataRd	 = 	 1'b0
;    2289		:	dataRd	 = 	 1'b0
;    2290		:	dataRd	 = 	 1'b0
;    2291		:	dataRd	 = 	 1'b0
;    2292		:	dataRd	 = 	 1'b1
;    2293		:	dataRd	 = 	 1'b0
;    2294		:	dataRd	 = 	 1'b0
;    2295		:	dataRd	 = 	 1'b0
;    2296		:	dataRd	 = 	 1'b0
;    2297		:	dataRd	 = 	 1'b0
;    2298		:	dataRd	 = 	 1'b0
;    2299		:	dataRd	 = 	 1'b0
;    2300		:	dataRd	 = 	 1'b0
;    2301		:	dataRd	 = 	 1'b0
;    2302		:	dataRd	 = 	 1'b0
;    2303		:	dataRd	 = 	 1'b0
;    2304		:	dataRd	 = 	 1'b0
;    2305		:	dataRd	 = 	 1'b0
;    2306		:	dataRd	 = 	 1'b0
;    2307		:	dataRd	 = 	 1'b0
;    2308		:	dataRd	 = 	 1'b1
;    2309		:	dataRd	 = 	 1'b0
;    2310		:	dataRd	 = 	 1'b0
;    2311		:	dataRd	 = 	 1'b0
;    2312		:	dataRd	 = 	 1'b0
;    2313		:	dataRd	 = 	 1'b0
;    2314		:	dataRd	 = 	 1'b0
;    2315		:	dataRd	 = 	 1'b0
;    2316		:	dataRd	 = 	 1'b0
;    2317		:	dataRd	 = 	 1'b0
;    2318		:	dataRd	 = 	 1'b0
;    2319		:	dataRd	 = 	 1'b0
;    2320		:	dataRd	 = 	 1'b0
;    2321		:	dataRd	 = 	 1'b0
;    2322		:	dataRd	 = 	 1'b0
;    2323		:	dataRd	 = 	 1'b0
;    2324		:	dataRd	 = 	 1'b1
;    2325		:	dataRd	 = 	 1'b0
;    2326		:	dataRd	 = 	 1'b0
;    2327		:	dataRd	 = 	 1'b0
;    2328		:	dataRd	 = 	 1'b0
;    2329		:	dataRd	 = 	 1'b0
;    2330		:	dataRd	 = 	 1'b0
;    2331		:	dataRd	 = 	 1'b0
;    2332		:	dataRd	 = 	 1'b0
;    2333		:	dataRd	 = 	 1'b0
;    2334		:	dataRd	 = 	 1'b0
;    2335		:	dataRd	 = 	 1'b0
;    2336		:	dataRd	 = 	 1'b0
;    2337		:	dataRd	 = 	 1'b0
;    2338		:	dataRd	 = 	 1'b0
;    2339		:	dataRd	 = 	 1'b0
;    2340		:	dataRd	 = 	 1'b1
;    2341		:	dataRd	 = 	 1'b0
;    2342		:	dataRd	 = 	 1'b0
;    2343		:	dataRd	 = 	 1'b0
;    2344		:	dataRd	 = 	 1'b0
;    2345		:	dataRd	 = 	 1'b0
;    2346		:	dataRd	 = 	 1'b0
;    2347		:	dataRd	 = 	 1'b0
;    2348		:	dataRd	 = 	 1'b0
;    2349		:	dataRd	 = 	 1'b0
;    2350		:	dataRd	 = 	 1'b0
;    2351		:	dataRd	 = 	 1'b0
;    2352		:	dataRd	 = 	 1'b0
;    2353		:	dataRd	 = 	 1'b0
;    2354		:	dataRd	 = 	 1'b0
;    2355		:	dataRd	 = 	 1'b0
;    2356		:	dataRd	 = 	 1'b1
;    2357		:	dataRd	 = 	 1'b0
;    2358		:	dataRd	 = 	 1'b0
;    2359		:	dataRd	 = 	 1'b0
;    2360		:	dataRd	 = 	 1'b0
;    2361		:	dataRd	 = 	 1'b0
;    2362		:	dataRd	 = 	 1'b0
;    2363		:	dataRd	 = 	 1'b0
;    2364		:	dataRd	 = 	 1'b0
;    2365		:	dataRd	 = 	 1'b0
;    2366		:	dataRd	 = 	 1'b0
;    2367		:	dataRd	 = 	 1'b0
;    2368		:	dataRd	 = 	 1'b0
;    2369		:	dataRd	 = 	 1'b0
;    2370		:	dataRd	 = 	 1'b0
;    2371		:	dataRd	 = 	 1'b0
;    2372		:	dataRd	 = 	 1'b1
;    2373		:	dataRd	 = 	 1'b0
;    2374		:	dataRd	 = 	 1'b0
;    2375		:	dataRd	 = 	 1'b0
;    2376		:	dataRd	 = 	 1'b0
;    2377		:	dataRd	 = 	 1'b0
;    2378		:	dataRd	 = 	 1'b0
;    2379		:	dataRd	 = 	 1'b0
;    2380		:	dataRd	 = 	 1'b0
;    2381		:	dataRd	 = 	 1'b0
;    2382		:	dataRd	 = 	 1'b0
;    2383		:	dataRd	 = 	 1'b0
;    2384		:	dataRd	 = 	 1'b0
;    2385		:	dataRd	 = 	 1'b0
;    2386		:	dataRd	 = 	 1'b0
;    2387		:	dataRd	 = 	 1'b0
;    2388		:	dataRd	 = 	 1'b1
;    2389		:	dataRd	 = 	 1'b0
;    2390		:	dataRd	 = 	 1'b0
;    2391		:	dataRd	 = 	 1'b0
;    2392		:	dataRd	 = 	 1'b0
;    2393		:	dataRd	 = 	 1'b0
;    2394		:	dataRd	 = 	 1'b0
;    2395		:	dataRd	 = 	 1'b0
;    2396		:	dataRd	 = 	 1'b0
;    2397		:	dataRd	 = 	 1'b0
;    2398		:	dataRd	 = 	 1'b0
;    2399		:	dataRd	 = 	 1'b0
;    2400		:	dataRd	 = 	 1'b0
;    2401		:	dataRd	 = 	 1'b0
;    2402		:	dataRd	 = 	 1'b0
;    2403		:	dataRd	 = 	 1'b0
;    2404		:	dataRd	 = 	 1'b1
;    2405		:	dataRd	 = 	 1'b0
;    2406		:	dataRd	 = 	 1'b0
;    2407		:	dataRd	 = 	 1'b0
;    2408		:	dataRd	 = 	 1'b0
;    2409		:	dataRd	 = 	 1'b0
;    2410		:	dataRd	 = 	 1'b0
;    2411		:	dataRd	 = 	 1'b0
;    2412		:	dataRd	 = 	 1'b0
;    2413		:	dataRd	 = 	 1'b0
;    2414		:	dataRd	 = 	 1'b0
;    2415		:	dataRd	 = 	 1'b0
;    2416		:	dataRd	 = 	 1'b0
;    2417		:	dataRd	 = 	 1'b0
;    2418		:	dataRd	 = 	 1'b0
;    2419		:	dataRd	 = 	 1'b0
;    2420		:	dataRd	 = 	 1'b1
;    2421		:	dataRd	 = 	 1'b0
;    2422		:	dataRd	 = 	 1'b0
;    2423		:	dataRd	 = 	 1'b0
;    2424		:	dataRd	 = 	 1'b0
;    2425		:	dataRd	 = 	 1'b0
;    2426		:	dataRd	 = 	 1'b0
;    2427		:	dataRd	 = 	 1'b0
;    2428		:	dataRd	 = 	 1'b0
;    2429		:	dataRd	 = 	 1'b0
;    2430		:	dataRd	 = 	 1'b0
;    2431		:	dataRd	 = 	 1'b0
;    2432		:	dataRd	 = 	 1'b0
;    2433		:	dataRd	 = 	 1'b0
;    2434		:	dataRd	 = 	 1'b0
;    2435		:	dataRd	 = 	 1'b0
;    2436		:	dataRd	 = 	 1'b1
;    2437		:	dataRd	 = 	 1'b0
;    2438		:	dataRd	 = 	 1'b0
;    2439		:	dataRd	 = 	 1'b0
;    2440		:	dataRd	 = 	 1'b0
;    2441		:	dataRd	 = 	 1'b0
;    2442		:	dataRd	 = 	 1'b0
;    2443		:	dataRd	 = 	 1'b0
;    2444		:	dataRd	 = 	 1'b0
;    2445		:	dataRd	 = 	 1'b0
;    2446		:	dataRd	 = 	 1'b0
;    2447		:	dataRd	 = 	 1'b0
;    2448		:	dataRd	 = 	 1'b0
;    2449		:	dataRd	 = 	 1'b0
;    2450		:	dataRd	 = 	 1'b0
;    2451		:	dataRd	 = 	 1'b0
;    2452		:	dataRd	 = 	 1'b1
;    2453		:	dataRd	 = 	 1'b0
;    2454		:	dataRd	 = 	 1'b0
;    2455		:	dataRd	 = 	 1'b0
;    2456		:	dataRd	 = 	 1'b0
;    2457		:	dataRd	 = 	 1'b0
;    2458		:	dataRd	 = 	 1'b0
;    2459		:	dataRd	 = 	 1'b0
;    2460		:	dataRd	 = 	 1'b0
;    2461		:	dataRd	 = 	 1'b0
;    2462		:	dataRd	 = 	 1'b0
;    2463		:	dataRd	 = 	 1'b0
;    2464		:	dataRd	 = 	 1'b0
;    2465		:	dataRd	 = 	 1'b0
;    2466		:	dataRd	 = 	 1'b0
;    2467		:	dataRd	 = 	 1'b0
;    2468		:	dataRd	 = 	 1'b1
;    2469		:	dataRd	 = 	 1'b0
;    2470		:	dataRd	 = 	 1'b0
;    2471		:	dataRd	 = 	 1'b0
;    2472		:	dataRd	 = 	 1'b0
;    2473		:	dataRd	 = 	 1'b0
;    2474		:	dataRd	 = 	 1'b0
;    2475		:	dataRd	 = 	 1'b0
;    2476		:	dataRd	 = 	 1'b0
;    2477		:	dataRd	 = 	 1'b0
;    2478		:	dataRd	 = 	 1'b0
;    2479		:	dataRd	 = 	 1'b0
;    2480		:	dataRd	 = 	 1'b0
;    2481		:	dataRd	 = 	 1'b0
;    2482		:	dataRd	 = 	 1'b0
;    2483		:	dataRd	 = 	 1'b0
;    2484		:	dataRd	 = 	 1'b1
;    2485		:	dataRd	 = 	 1'b0
;    2486		:	dataRd	 = 	 1'b0
;    2487		:	dataRd	 = 	 1'b0
;    2488		:	dataRd	 = 	 1'b0
;    2489		:	dataRd	 = 	 1'b0
;    2490		:	dataRd	 = 	 1'b0
;    2491		:	dataRd	 = 	 1'b0
;    2492		:	dataRd	 = 	 1'b0
;    2493		:	dataRd	 = 	 1'b0
;    2494		:	dataRd	 = 	 1'b0
;    2495		:	dataRd	 = 	 1'b0
;    2496		:	dataRd	 = 	 1'b0
;    2497		:	dataRd	 = 	 1'b0
;    2498		:	dataRd	 = 	 1'b0
;    2499		:	dataRd	 = 	 1'b0
;    2500		:	dataRd	 = 	 1'b1
;    2501		:	dataRd	 = 	 1'b0
;    2502		:	dataRd	 = 	 1'b0
;    2503		:	dataRd	 = 	 1'b0
;    2504		:	dataRd	 = 	 1'b0
;    2505		:	dataRd	 = 	 1'b0
;    2506		:	dataRd	 = 	 1'b0
;    2507		:	dataRd	 = 	 1'b0
;    2508		:	dataRd	 = 	 1'b0
;    2509		:	dataRd	 = 	 1'b0
;    2510		:	dataRd	 = 	 1'b0
;    2511		:	dataRd	 = 	 1'b0
;    2512		:	dataRd	 = 	 1'b0
;    2513		:	dataRd	 = 	 1'b0
;    2514		:	dataRd	 = 	 1'b0
;    2515		:	dataRd	 = 	 1'b0
;    2516		:	dataRd	 = 	 1'b1
;    2517		:	dataRd	 = 	 1'b0
;    2518		:	dataRd	 = 	 1'b0
;    2519		:	dataRd	 = 	 1'b0
;    2520		:	dataRd	 = 	 1'b0
;    2521		:	dataRd	 = 	 1'b0
;    2522		:	dataRd	 = 	 1'b0
;    2523		:	dataRd	 = 	 1'b0
;    2524		:	dataRd	 = 	 1'b0
;    2525		:	dataRd	 = 	 1'b0
;    2526		:	dataRd	 = 	 1'b0
;    2527		:	dataRd	 = 	 1'b0
;    2528		:	dataRd	 = 	 1'b0
;    2529		:	dataRd	 = 	 1'b0
;    2530		:	dataRd	 = 	 1'b0
;    2531		:	dataRd	 = 	 1'b0
;    2532		:	dataRd	 = 	 1'b1
;    2533		:	dataRd	 = 	 1'b0
;    2534		:	dataRd	 = 	 1'b0
;    2535		:	dataRd	 = 	 1'b0
;    2536		:	dataRd	 = 	 1'b0
;    2537		:	dataRd	 = 	 1'b0
;    2538		:	dataRd	 = 	 1'b0
;    2539		:	dataRd	 = 	 1'b0
;    2540		:	dataRd	 = 	 1'b0
;    2541		:	dataRd	 = 	 1'b0
;    2542		:	dataRd	 = 	 1'b0
;    2543		:	dataRd	 = 	 1'b0
;    2544		:	dataRd	 = 	 1'b0
;    2545		:	dataRd	 = 	 1'b0
;    2546		:	dataRd	 = 	 1'b0
;    2547		:	dataRd	 = 	 1'b0
;    2548		:	dataRd	 = 	 1'b1
;    2549		:	dataRd	 = 	 1'b0
;    2550		:	dataRd	 = 	 1'b0
;    2551		:	dataRd	 = 	 1'b0
;    2552		:	dataRd	 = 	 1'b0
;    2553		:	dataRd	 = 	 1'b0
;    2554		:	dataRd	 = 	 1'b0
;    2555		:	dataRd	 = 	 1'b0
;    2556		:	dataRd	 = 	 1'b0
;    2557		:	dataRd	 = 	 1'b0
;    2558		:	dataRd	 = 	 1'b0
;    2559		:	dataRd	 = 	 1'b0
;    2560		:	dataRd	 = 	 1'b0
;    2561		:	dataRd	 = 	 1'b0
;    2562		:	dataRd	 = 	 1'b0
;    2563		:	dataRd	 = 	 1'b0
;    2564		:	dataRd	 = 	 1'b1
;    2565		:	dataRd	 = 	 1'b0
;    2566		:	dataRd	 = 	 1'b0
;    2567		:	dataRd	 = 	 1'b0
;    2568		:	dataRd	 = 	 1'b0
;    2569		:	dataRd	 = 	 1'b0
;    2570		:	dataRd	 = 	 1'b0
;    2571		:	dataRd	 = 	 1'b0
;    2572		:	dataRd	 = 	 1'b0
;    2573		:	dataRd	 = 	 1'b0
;    2574		:	dataRd	 = 	 1'b0
;    2575		:	dataRd	 = 	 1'b0
;    2576		:	dataRd	 = 	 1'b0
;    2577		:	dataRd	 = 	 1'b0
;    2578		:	dataRd	 = 	 1'b0
;    2579		:	dataRd	 = 	 1'b0
;    2580		:	dataRd	 = 	 1'b1
;    2581		:	dataRd	 = 	 1'b0
;    2582		:	dataRd	 = 	 1'b0
;    2583		:	dataRd	 = 	 1'b0
;    2584		:	dataRd	 = 	 1'b0
;    2585		:	dataRd	 = 	 1'b0
;    2586		:	dataRd	 = 	 1'b0
;    2587		:	dataRd	 = 	 1'b0
;    2588		:	dataRd	 = 	 1'b0
;    2589		:	dataRd	 = 	 1'b0
;    2590		:	dataRd	 = 	 1'b0
;    2591		:	dataRd	 = 	 1'b0
;    2592		:	dataRd	 = 	 1'b0
;    2593		:	dataRd	 = 	 1'b0
;    2594		:	dataRd	 = 	 1'b0
;    2595		:	dataRd	 = 	 1'b0
;    2596		:	dataRd	 = 	 1'b1
;    2597		:	dataRd	 = 	 1'b0
;    2598		:	dataRd	 = 	 1'b0
;    2599		:	dataRd	 = 	 1'b0
;    2600		:	dataRd	 = 	 1'b0
;    2601		:	dataRd	 = 	 1'b0
;    2602		:	dataRd	 = 	 1'b0
;    2603		:	dataRd	 = 	 1'b0
;    2604		:	dataRd	 = 	 1'b0
;    2605		:	dataRd	 = 	 1'b0
;    2606		:	dataRd	 = 	 1'b0
;    2607		:	dataRd	 = 	 1'b0
;    2608		:	dataRd	 = 	 1'b0
;    2609		:	dataRd	 = 	 1'b0
;    2610		:	dataRd	 = 	 1'b0
;    2611		:	dataRd	 = 	 1'b0
;    2612		:	dataRd	 = 	 1'b1
;    2613		:	dataRd	 = 	 1'b0
;    2614		:	dataRd	 = 	 1'b0
;    2615		:	dataRd	 = 	 1'b0
;    2616		:	dataRd	 = 	 1'b0
;    2617		:	dataRd	 = 	 1'b0
;    2618		:	dataRd	 = 	 1'b0
;    2619		:	dataRd	 = 	 1'b0
;    2620		:	dataRd	 = 	 1'b0
;    2621		:	dataRd	 = 	 1'b0
;    2622		:	dataRd	 = 	 1'b0
;    2623		:	dataRd	 = 	 1'b0
;    2624		:	dataRd	 = 	 1'b0
;    2625		:	dataRd	 = 	 1'b0
;    2626		:	dataRd	 = 	 1'b0
;    2627		:	dataRd	 = 	 1'b0
;    2628		:	dataRd	 = 	 1'b1
;    2629		:	dataRd	 = 	 1'b0
;    2630		:	dataRd	 = 	 1'b0
;    2631		:	dataRd	 = 	 1'b0
;    2632		:	dataRd	 = 	 1'b0
;    2633		:	dataRd	 = 	 1'b0
;    2634		:	dataRd	 = 	 1'b0
;    2635		:	dataRd	 = 	 1'b0
;    2636		:	dataRd	 = 	 1'b0
;    2637		:	dataRd	 = 	 1'b0
;    2638		:	dataRd	 = 	 1'b0
;    2639		:	dataRd	 = 	 1'b0
;    2640		:	dataRd	 = 	 1'b0
;    2641		:	dataRd	 = 	 1'b0
;    2642		:	dataRd	 = 	 1'b0
;    2643		:	dataRd	 = 	 1'b0
;    2644		:	dataRd	 = 	 1'b1
;    2645		:	dataRd	 = 	 1'b0
;    2646		:	dataRd	 = 	 1'b0
;    2647		:	dataRd	 = 	 1'b0
;    2648		:	dataRd	 = 	 1'b0
;    2649		:	dataRd	 = 	 1'b0
;    2650		:	dataRd	 = 	 1'b0
;    2651		:	dataRd	 = 	 1'b0
;    2652		:	dataRd	 = 	 1'b0
;    2653		:	dataRd	 = 	 1'b0
;    2654		:	dataRd	 = 	 1'b0
;    2655		:	dataRd	 = 	 1'b0
;    2656		:	dataRd	 = 	 1'b0
;    2657		:	dataRd	 = 	 1'b0
;    2658		:	dataRd	 = 	 1'b0
;    2659		:	dataRd	 = 	 1'b0
;    2660		:	dataRd	 = 	 1'b1
;    2661		:	dataRd	 = 	 1'b0
;    2662		:	dataRd	 = 	 1'b0
;    2663		:	dataRd	 = 	 1'b0
;    2664		:	dataRd	 = 	 1'b0
;    2665		:	dataRd	 = 	 1'b0
;    2666		:	dataRd	 = 	 1'b0
;    2667		:	dataRd	 = 	 1'b0
;    2668		:	dataRd	 = 	 1'b0
;    2669		:	dataRd	 = 	 1'b0
;    2670		:	dataRd	 = 	 1'b0
;    2671		:	dataRd	 = 	 1'b0
;    2672		:	dataRd	 = 	 1'b0
;    2673		:	dataRd	 = 	 1'b0
;    2674		:	dataRd	 = 	 1'b0
;    2675		:	dataRd	 = 	 1'b0
;    2676		:	dataRd	 = 	 1'b1
;    2677		:	dataRd	 = 	 1'b0
;    2678		:	dataRd	 = 	 1'b0
;    2679		:	dataRd	 = 	 1'b0
;    2680		:	dataRd	 = 	 1'b0
;    2681		:	dataRd	 = 	 1'b0
;    2682		:	dataRd	 = 	 1'b0
;    2683		:	dataRd	 = 	 1'b0
;    2684		:	dataRd	 = 	 1'b0
;    2685		:	dataRd	 = 	 1'b0
;    2686		:	dataRd	 = 	 1'b0
;    2687		:	dataRd	 = 	 1'b0
;    2688		:	dataRd	 = 	 1'b0
;    2689		:	dataRd	 = 	 1'b0
;    2690		:	dataRd	 = 	 1'b0
;    2691		:	dataRd	 = 	 1'b0
;    2692		:	dataRd	 = 	 1'b1
;    2693		:	dataRd	 = 	 1'b0
;    2694		:	dataRd	 = 	 1'b0
;    2695		:	dataRd	 = 	 1'b0
;    2696		:	dataRd	 = 	 1'b0
;    2697		:	dataRd	 = 	 1'b0
;    2698		:	dataRd	 = 	 1'b0
;    2699		:	dataRd	 = 	 1'b0
;    2700		:	dataRd	 = 	 1'b0
;    2701		:	dataRd	 = 	 1'b0
;    2702		:	dataRd	 = 	 1'b0
;    2703		:	dataRd	 = 	 1'b0
;    2704		:	dataRd	 = 	 1'b0
;    2705		:	dataRd	 = 	 1'b0
;    2706		:	dataRd	 = 	 1'b0
;    2707		:	dataRd	 = 	 1'b0
;    2708		:	dataRd	 = 	 1'b1
;    2709		:	dataRd	 = 	 1'b0
;    2710		:	dataRd	 = 	 1'b0
;    2711		:	dataRd	 = 	 1'b0
;    2712		:	dataRd	 = 	 1'b0
;    2713		:	dataRd	 = 	 1'b0
;    2714		:	dataRd	 = 	 1'b0
;    2715		:	dataRd	 = 	 1'b0
;    2716		:	dataRd	 = 	 1'b0
;    2717		:	dataRd	 = 	 1'b0
;    2718		:	dataRd	 = 	 1'b0
;    2719		:	dataRd	 = 	 1'b0
;    2720		:	dataRd	 = 	 1'b0
;    2721		:	dataRd	 = 	 1'b0
;    2722		:	dataRd	 = 	 1'b0
;    2723		:	dataRd	 = 	 1'b0
;    2724		:	dataRd	 = 	 1'b0
;    2725		:	dataRd	 = 	 1'b0
;    2726		:	dataRd	 = 	 1'b0
;    2727		:	dataRd	 = 	 1'b0
;    2728		:	dataRd	 = 	 1'b0
;    2729		:	dataRd	 = 	 1'b0
;    2730		:	dataRd	 = 	 1'b0
;    2731		:	dataRd	 = 	 1'b0
;    2732		:	dataRd	 = 	 1'b0
;    2733		:	dataRd	 = 	 1'b0
;    2734		:	dataRd	 = 	 1'b0
;    2735		:	dataRd	 = 	 1'b0
;    2736		:	dataRd	 = 	 1'b0
;    2737		:	dataRd	 = 	 1'b0
;    2738		:	dataRd	 = 	 1'b0
;    2739		:	dataRd	 = 	 1'b0
;    2740		:	dataRd	 = 	 1'b0
;    2741		:	dataRd	 = 	 1'b0
;    2742		:	dataRd	 = 	 1'b0
;    2743		:	dataRd	 = 	 1'b0
;    2744		:	dataRd	 = 	 1'b0
;    2745		:	dataRd	 = 	 1'b0
;    2746		:	dataRd	 = 	 1'b0
;    2747		:	dataRd	 = 	 1'b0
;    2748		:	dataRd	 = 	 1'b0
;    2749		:	dataRd	 = 	 1'b0
;    2750		:	dataRd	 = 	 1'b0
;    2751		:	dataRd	 = 	 1'b0
;    2752		:	dataRd	 = 	 1'b0
;    2753		:	dataRd	 = 	 1'b0
;    2754		:	dataRd	 = 	 1'b0
;    2755		:	dataRd	 = 	 1'b0
;    2756		:	dataRd	 = 	 1'b0
;    2757		:	dataRd	 = 	 1'b0
;    2758		:	dataRd	 = 	 1'b0
;    2759		:	dataRd	 = 	 1'b0
;    2760		:	dataRd	 = 	 1'b0
;    2761		:	dataRd	 = 	 1'b0
;    2762		:	dataRd	 = 	 1'b0
;    2763		:	dataRd	 = 	 1'b0
;    2764		:	dataRd	 = 	 1'b0
;    2765		:	dataRd	 = 	 1'b0
;    2766		:	dataRd	 = 	 1'b0
;    2767		:	dataRd	 = 	 1'b0
;    2768		:	dataRd	 = 	 1'b0
;    2769		:	dataRd	 = 	 1'b0
;    2770		:	dataRd	 = 	 1'b0
;    2771		:	dataRd	 = 	 1'b0
;    2772		:	dataRd	 = 	 1'b0
;    2773		:	dataRd	 = 	 1'b0
;    2774		:	dataRd	 = 	 1'b0
;    2775		:	dataRd	 = 	 1'b1
;    2776		:	dataRd	 = 	 1'b0
;    2777		:	dataRd	 = 	 1'b0
;    2778		:	dataRd	 = 	 1'b0
;    2779		:	dataRd	 = 	 1'b0
;    2780		:	dataRd	 = 	 1'b0
;    2781		:	dataRd	 = 	 1'b0
;    2782		:	dataRd	 = 	 1'b0
;    2783		:	dataRd	 = 	 1'b0
;    2784		:	dataRd	 = 	 1'b0
;    2785		:	dataRd	 = 	 1'b0
;    2786		:	dataRd	 = 	 1'b0
;    2787		:	dataRd	 = 	 1'b0
;    2788		:	dataRd	 = 	 1'b0
;    2789		:	dataRd	 = 	 1'b0
;    2790		:	dataRd	 = 	 1'b0
;    2791		:	dataRd	 = 	 1'b0
;    2792		:	dataRd	 = 	 1'b0
;    2793		:	dataRd	 = 	 1'b0
;    2794		:	dataRd	 = 	 1'b0
;    2795		:	dataRd	 = 	 1'b0
;    2796		:	dataRd	 = 	 1'b0
;    2797		:	dataRd	 = 	 1'b0
;    2798		:	dataRd	 = 	 1'b0
;    2799		:	dataRd	 = 	 1'b0
;    2800		:	dataRd	 = 	 1'b0
;    2801		:	dataRd	 = 	 1'b0
;    2802		:	dataRd	 = 	 1'b0
;    2803		:	dataRd	 = 	 1'b0
;    2804		:	dataRd	 = 	 1'b0
;    2805		:	dataRd	 = 	 1'b0
;    2806		:	dataRd	 = 	 1'b0
;    2807		:	dataRd	 = 	 1'b0
;    2808		:	dataRd	 = 	 1'b0
;    2809		:	dataRd	 = 	 1'b0
;    2810		:	dataRd	 = 	 1'b0
;    2811		:	dataRd	 = 	 1'b0
;    2812		:	dataRd	 = 	 1'b0
;    2813		:	dataRd	 = 	 1'b0
;    2814		:	dataRd	 = 	 1'b0
;    2815		:	dataRd	 = 	 1'b0
;    2816		:	dataRd	 = 	 1'b0
;    2817		:	dataRd	 = 	 1'b0
;    2818		:	dataRd	 = 	 1'b0
;    2819		:	dataRd	 = 	 1'b0
;    2820		:	dataRd	 = 	 1'b0
;    2821		:	dataRd	 = 	 1'b0
;    2822		:	dataRd	 = 	 1'b0
;    2823		:	dataRd	 = 	 1'b0
;    2824		:	dataRd	 = 	 1'b0
;    2825		:	dataRd	 = 	 1'b0
;    2826		:	dataRd	 = 	 1'b0
;    2827		:	dataRd	 = 	 1'b0
;    2828		:	dataRd	 = 	 1'b0
;    2829		:	dataRd	 = 	 1'b0
;    2830		:	dataRd	 = 	 1'b0
;    2831		:	dataRd	 = 	 1'b0
;    2832		:	dataRd	 = 	 1'b0
;    2833		:	dataRd	 = 	 1'b0
;    2834		:	dataRd	 = 	 1'b0
;    2835		:	dataRd	 = 	 1'b0
;    2836		:	dataRd	 = 	 1'b0
;    2837		:	dataRd	 = 	 1'b0
;    2838		:	dataRd	 = 	 1'b0
;    2839		:	dataRd	 = 	 1'b0
;    2840		:	dataRd	 = 	 1'b0
;    2841		:	dataRd	 = 	 1'b0
;    2842		:	dataRd	 = 	 1'b1
;    2843		:	dataRd	 = 	 1'b0
;    2844		:	dataRd	 = 	 1'b0
;    2845		:	dataRd	 = 	 1'b0
;    2846		:	dataRd	 = 	 1'b0
;    2847		:	dataRd	 = 	 1'b0
;    2848		:	dataRd	 = 	 1'b0
;    2849		:	dataRd	 = 	 1'b0
;    2850		:	dataRd	 = 	 1'b0
;    2851		:	dataRd	 = 	 1'b0
;    2852		:	dataRd	 = 	 1'b0
;    2853		:	dataRd	 = 	 1'b0
;    2854		:	dataRd	 = 	 1'b0
;    2855		:	dataRd	 = 	 1'b0
;    2856		:	dataRd	 = 	 1'b0
;    2857		:	dataRd	 = 	 1'b0
;    2858		:	dataRd	 = 	 1'b0
;    2859		:	dataRd	 = 	 1'b0
;    2860		:	dataRd	 = 	 1'b0
;    2861		:	dataRd	 = 	 1'b0
;    2862		:	dataRd	 = 	 1'b0
;    2863		:	dataRd	 = 	 1'b0
;    2864		:	dataRd	 = 	 1'b0
;    2865		:	dataRd	 = 	 1'b0
;    2866		:	dataRd	 = 	 1'b0
;    2867		:	dataRd	 = 	 1'b0
;    2868		:	dataRd	 = 	 1'b0
;    2869		:	dataRd	 = 	 1'b0
;    2870		:	dataRd	 = 	 1'b0
;    2871		:	dataRd	 = 	 1'b0
;    2872		:	dataRd	 = 	 1'b0
;    2873		:	dataRd	 = 	 1'b0
;    2874		:	dataRd	 = 	 1'b0
;    2875		:	dataRd	 = 	 1'b0
;    2876		:	dataRd	 = 	 1'b0
;    2877		:	dataRd	 = 	 1'b0
;    2878		:	dataRd	 = 	 1'b0
;    2879		:	dataRd	 = 	 1'b0
;    2880		:	dataRd	 = 	 1'b0
;    2881		:	dataRd	 = 	 1'b0
;    2882		:	dataRd	 = 	 1'b0
;    2883		:	dataRd	 = 	 1'b0
;    2884		:	dataRd	 = 	 1'b0
;    2885		:	dataRd	 = 	 1'b0
;    2886		:	dataRd	 = 	 1'b0
;    2887		:	dataRd	 = 	 1'b0
;    2888		:	dataRd	 = 	 1'b0
;    2889		:	dataRd	 = 	 1'b0
;    2890		:	dataRd	 = 	 1'b0
;    2891		:	dataRd	 = 	 1'b0
;    2892		:	dataRd	 = 	 1'b0
;    2893		:	dataRd	 = 	 1'b0
;    2894		:	dataRd	 = 	 1'b0
;    2895		:	dataRd	 = 	 1'b0
;    2896		:	dataRd	 = 	 1'b0
;    2897		:	dataRd	 = 	 1'b0
;    2898		:	dataRd	 = 	 1'b0
;    2899		:	dataRd	 = 	 1'b0
;    2900		:	dataRd	 = 	 1'b0
;    2901		:	dataRd	 = 	 1'b0
;    2902		:	dataRd	 = 	 1'b0
;    2903		:	dataRd	 = 	 1'b0
;    2904		:	dataRd	 = 	 1'b0
;    2905		:	dataRd	 = 	 1'b0
;    2906		:	dataRd	 = 	 1'b0
;    2907		:	dataRd	 = 	 1'b0
;    2908		:	dataRd	 = 	 1'b0
;    2909		:	dataRd	 = 	 1'b1
;    2910		:	dataRd	 = 	 1'b0
;    2911		:	dataRd	 = 	 1'b0
;    2912		:	dataRd	 = 	 1'b0
;    2913		:	dataRd	 = 	 1'b0
;    2914		:	dataRd	 = 	 1'b0
;    2915		:	dataRd	 = 	 1'b0
;    2916		:	dataRd	 = 	 1'b0
;    2917		:	dataRd	 = 	 1'b0
;    2918		:	dataRd	 = 	 1'b0
;    2919		:	dataRd	 = 	 1'b0
;    2920		:	dataRd	 = 	 1'b0
;    2921		:	dataRd	 = 	 1'b0
;    2922		:	dataRd	 = 	 1'b0
;    2923		:	dataRd	 = 	 1'b0
;    2924		:	dataRd	 = 	 1'b0
;    2925		:	dataRd	 = 	 1'b0
;    2926		:	dataRd	 = 	 1'b0
;    2927		:	dataRd	 = 	 1'b0
;    2928		:	dataRd	 = 	 1'b0
;    2929		:	dataRd	 = 	 1'b0
;    2930		:	dataRd	 = 	 1'b0
;    2931		:	dataRd	 = 	 1'b0
;    2932		:	dataRd	 = 	 1'b0
;    2933		:	dataRd	 = 	 1'b0
;    2934		:	dataRd	 = 	 1'b0
;    2935		:	dataRd	 = 	 1'b0
;    2936		:	dataRd	 = 	 1'b0
;    2937		:	dataRd	 = 	 1'b0
;    2938		:	dataRd	 = 	 1'b0
;    2939		:	dataRd	 = 	 1'b0
;    2940		:	dataRd	 = 	 1'b0
;    2941		:	dataRd	 = 	 1'b0
;    2942		:	dataRd	 = 	 1'b0
;    2943		:	dataRd	 = 	 1'b0
;    2944		:	dataRd	 = 	 1'b0
;    2945		:	dataRd	 = 	 1'b0
;    2946		:	dataRd	 = 	 1'b0
;    2947		:	dataRd	 = 	 1'b0
;    2948		:	dataRd	 = 	 1'b0
;    2949		:	dataRd	 = 	 1'b0
;    2950		:	dataRd	 = 	 1'b0
;    2951		:	dataRd	 = 	 1'b0
;    2952		:	dataRd	 = 	 1'b0
;    2953		:	dataRd	 = 	 1'b0
;    2954		:	dataRd	 = 	 1'b0
;    2955		:	dataRd	 = 	 1'b0
;    2956		:	dataRd	 = 	 1'b0
;    2957		:	dataRd	 = 	 1'b0
;    2958		:	dataRd	 = 	 1'b0
;    2959		:	dataRd	 = 	 1'b0
;    2960		:	dataRd	 = 	 1'b0
;    2961		:	dataRd	 = 	 1'b0
;    2962		:	dataRd	 = 	 1'b0
;    2963		:	dataRd	 = 	 1'b0
;    2964		:	dataRd	 = 	 1'b0
;    2965		:	dataRd	 = 	 1'b0
;    2966		:	dataRd	 = 	 1'b0
;    2967		:	dataRd	 = 	 1'b0
;    2968		:	dataRd	 = 	 1'b0
;    2969		:	dataRd	 = 	 1'b0
;    2970		:	dataRd	 = 	 1'b0
;    2971		:	dataRd	 = 	 1'b0
;    2972		:	dataRd	 = 	 1'b0
;    2973		:	dataRd	 = 	 1'b0
;    2974		:	dataRd	 = 	 1'b0
;    2975		:	dataRd	 = 	 1'b0
;    2976		:	dataRd	 = 	 1'b1
;    2977		:	dataRd	 = 	 1'b0
;    2978		:	dataRd	 = 	 1'b0
;    2979		:	dataRd	 = 	 1'b0
;    2980		:	dataRd	 = 	 1'b0
;    2981		:	dataRd	 = 	 1'b0
;    2982		:	dataRd	 = 	 1'b0
;    2983		:	dataRd	 = 	 1'b0
;    2984		:	dataRd	 = 	 1'b0
;    2985		:	dataRd	 = 	 1'b0
;    2986		:	dataRd	 = 	 1'b0
;    2987		:	dataRd	 = 	 1'b0
;    2988		:	dataRd	 = 	 1'b0
;    2989		:	dataRd	 = 	 1'b0
;    2990		:	dataRd	 = 	 1'b0
;    2991		:	dataRd	 = 	 1'b0
;    2992		:	dataRd	 = 	 1'b0
;    2993		:	dataRd	 = 	 1'b0
;    2994		:	dataRd	 = 	 1'b0
;    2995		:	dataRd	 = 	 1'b0
;    2996		:	dataRd	 = 	 1'b0
;    2997		:	dataRd	 = 	 1'b0
;    2998		:	dataRd	 = 	 1'b0
;    2999		:	dataRd	 = 	 1'b0
;    3000		:	dataRd	 = 	 1'b0
;    3001		:	dataRd	 = 	 1'b0
;    3002		:	dataRd	 = 	 1'b0
;    3003		:	dataRd	 = 	 1'b0
;    3004		:	dataRd	 = 	 1'b0
;    3005		:	dataRd	 = 	 1'b0
;    3006		:	dataRd	 = 	 1'b0
;    3007		:	dataRd	 = 	 1'b0
;    3008		:	dataRd	 = 	 1'b0
;    3009		:	dataRd	 = 	 1'b0
;    3010		:	dataRd	 = 	 1'b0
;    3011		:	dataRd	 = 	 1'b0
;    3012		:	dataRd	 = 	 1'b0
;    3013		:	dataRd	 = 	 1'b0
;    3014		:	dataRd	 = 	 1'b0
;    3015		:	dataRd	 = 	 1'b0
;    3016		:	dataRd	 = 	 1'b0
;    3017		:	dataRd	 = 	 1'b0
;    3018		:	dataRd	 = 	 1'b0
;    3019		:	dataRd	 = 	 1'b0
;    3020		:	dataRd	 = 	 1'b0
;    3021		:	dataRd	 = 	 1'b0
;    3022		:	dataRd	 = 	 1'b0
;    3023		:	dataRd	 = 	 1'b0
;    3024		:	dataRd	 = 	 1'b0
;    3025		:	dataRd	 = 	 1'b0
;    3026		:	dataRd	 = 	 1'b0
;    3027		:	dataRd	 = 	 1'b0
;    3028		:	dataRd	 = 	 1'b0
;    3029		:	dataRd	 = 	 1'b0
;    3030		:	dataRd	 = 	 1'b0
;    3031		:	dataRd	 = 	 1'b0
;    3032		:	dataRd	 = 	 1'b0
;    3033		:	dataRd	 = 	 1'b0
;    3034		:	dataRd	 = 	 1'b0
;    3035		:	dataRd	 = 	 1'b0
;    3036		:	dataRd	 = 	 1'b0
;    3037		:	dataRd	 = 	 1'b0
;    3038		:	dataRd	 = 	 1'b0
;    3039		:	dataRd	 = 	 1'b0
;    3040		:	dataRd	 = 	 1'b0
;    3041		:	dataRd	 = 	 1'b0
;    3042		:	dataRd	 = 	 1'b0
;    3043		:	dataRd	 = 	 1'b1
;    3044		:	dataRd	 = 	 1'b0
;    3045		:	dataRd	 = 	 1'b0
;    3046		:	dataRd	 = 	 1'b0
;    3047		:	dataRd	 = 	 1'b0
;    3048		:	dataRd	 = 	 1'b0
;    3049		:	dataRd	 = 	 1'b0
;    3050		:	dataRd	 = 	 1'b0
;    3051		:	dataRd	 = 	 1'b0
;    3052		:	dataRd	 = 	 1'b0
;    3053		:	dataRd	 = 	 1'b0
;    3054		:	dataRd	 = 	 1'b0
;    3055		:	dataRd	 = 	 1'b0
;    3056		:	dataRd	 = 	 1'b0
;    3057		:	dataRd	 = 	 1'b0
;    3058		:	dataRd	 = 	 1'b0
;    3059		:	dataRd	 = 	 1'b0
;    3060		:	dataRd	 = 	 1'b0
;    3061		:	dataRd	 = 	 1'b0
;    3062		:	dataRd	 = 	 1'b0
;    3063		:	dataRd	 = 	 1'b0
;    3064		:	dataRd	 = 	 1'b0
;    3065		:	dataRd	 = 	 1'b0
;    3066		:	dataRd	 = 	 1'b0
;    3067		:	dataRd	 = 	 1'b0
;    3068		:	dataRd	 = 	 1'b0
;    3069		:	dataRd	 = 	 1'b0
;    3070		:	dataRd	 = 	 1'b0
;    3071		:	dataRd	 = 	 1'b0
;    3072		:	dataRd	 = 	 1'b0
;    3073		:	dataRd	 = 	 1'b0
;    3074		:	dataRd	 = 	 1'b0
;    3075		:	dataRd	 = 	 1'b0
;    3076		:	dataRd	 = 	 1'b0
;    3077		:	dataRd	 = 	 1'b0
;    3078		:	dataRd	 = 	 1'b0
;    3079		:	dataRd	 = 	 1'b0
;    3080		:	dataRd	 = 	 1'b0
;    3081		:	dataRd	 = 	 1'b0
;    3082		:	dataRd	 = 	 1'b0
;    3083		:	dataRd	 = 	 1'b0
;    3084		:	dataRd	 = 	 1'b0
;    3085		:	dataRd	 = 	 1'b0
;    3086		:	dataRd	 = 	 1'b0
;    3087		:	dataRd	 = 	 1'b0
;    3088		:	dataRd	 = 	 1'b0
;    3089		:	dataRd	 = 	 1'b0
;    3090		:	dataRd	 = 	 1'b0
;    3091		:	dataRd	 = 	 1'b0
;    3092		:	dataRd	 = 	 1'b0
;    3093		:	dataRd	 = 	 1'b0
;    3094		:	dataRd	 = 	 1'b0
;    3095		:	dataRd	 = 	 1'b0
;    3096		:	dataRd	 = 	 1'b0
;    3097		:	dataRd	 = 	 1'b0
;    3098		:	dataRd	 = 	 1'b0
;    3099		:	dataRd	 = 	 1'b0
;    3100		:	dataRd	 = 	 1'b0
;    3101		:	dataRd	 = 	 1'b0
;    3102		:	dataRd	 = 	 1'b0
;    3103		:	dataRd	 = 	 1'b0
;    3104		:	dataRd	 = 	 1'b0
;    3105		:	dataRd	 = 	 1'b0
;    3106		:	dataRd	 = 	 1'b0
;    3107		:	dataRd	 = 	 1'b0
;    3108		:	dataRd	 = 	 1'b0
;    3109		:	dataRd	 = 	 1'b0
;    3110		:	dataRd	 = 	 1'b1
;    3111		:	dataRd	 = 	 1'b0
;    3112		:	dataRd	 = 	 1'b0
;    3113		:	dataRd	 = 	 1'b0
;    3114		:	dataRd	 = 	 1'b0
;    3115		:	dataRd	 = 	 1'b0
;    3116		:	dataRd	 = 	 1'b0
;    3117		:	dataRd	 = 	 1'b0
;    3118		:	dataRd	 = 	 1'b0
;    3119		:	dataRd	 = 	 1'b0
;    3120		:	dataRd	 = 	 1'b0
;    3121		:	dataRd	 = 	 1'b0
;    3122		:	dataRd	 = 	 1'b0
;    3123		:	dataRd	 = 	 1'b0
;    3124		:	dataRd	 = 	 1'b0
;    3125		:	dataRd	 = 	 1'b0
;    3126		:	dataRd	 = 	 1'b0
;    3127		:	dataRd	 = 	 1'b0
;    3128		:	dataRd	 = 	 1'b0
;    3129		:	dataRd	 = 	 1'b0
;    3130		:	dataRd	 = 	 1'b0
;    3131		:	dataRd	 = 	 1'b0
;    3132		:	dataRd	 = 	 1'b0
;    3133		:	dataRd	 = 	 1'b0
;    3134		:	dataRd	 = 	 1'b0
;    3135		:	dataRd	 = 	 1'b0
;    3136		:	dataRd	 = 	 1'b0
;    3137		:	dataRd	 = 	 1'b0
;    3138		:	dataRd	 = 	 1'b0
;    3139		:	dataRd	 = 	 1'b0
;    3140		:	dataRd	 = 	 1'b0
;    3141		:	dataRd	 = 	 1'b0
;    3142		:	dataRd	 = 	 1'b0
;    3143		:	dataRd	 = 	 1'b0
;    3144		:	dataRd	 = 	 1'b0
;    3145		:	dataRd	 = 	 1'b0
;    3146		:	dataRd	 = 	 1'b0
;    3147		:	dataRd	 = 	 1'b0
;    3148		:	dataRd	 = 	 1'b0
;    3149		:	dataRd	 = 	 1'b0
;    3150		:	dataRd	 = 	 1'b0
;    3151		:	dataRd	 = 	 1'b0
;    3152		:	dataRd	 = 	 1'b0
;    3153		:	dataRd	 = 	 1'b0
;    3154		:	dataRd	 = 	 1'b0
;    3155		:	dataRd	 = 	 1'b0
;    3156		:	dataRd	 = 	 1'b0
;    3157		:	dataRd	 = 	 1'b0
;    3158		:	dataRd	 = 	 1'b0
;    3159		:	dataRd	 = 	 1'b0
;    3160		:	dataRd	 = 	 1'b0
;    3161		:	dataRd	 = 	 1'b0
;    3162		:	dataRd	 = 	 1'b0
;    3163		:	dataRd	 = 	 1'b0
;    3164		:	dataRd	 = 	 1'b0
;    3165		:	dataRd	 = 	 1'b0
;    3166		:	dataRd	 = 	 1'b0
;    3167		:	dataRd	 = 	 1'b0
;    3168		:	dataRd	 = 	 1'b0
;    3169		:	dataRd	 = 	 1'b0
;    3170		:	dataRd	 = 	 1'b0
;    3171		:	dataRd	 = 	 1'b0
;    3172		:	dataRd	 = 	 1'b0
;    3173		:	dataRd	 = 	 1'b0
;    3174		:	dataRd	 = 	 1'b0
;    3175		:	dataRd	 = 	 1'b0
;    3176		:	dataRd	 = 	 1'b0
;    3177		:	dataRd	 = 	 1'b1
;    3178		:	dataRd	 = 	 1'b0
;    3179		:	dataRd	 = 	 1'b0
;    3180		:	dataRd	 = 	 1'b0
;    3181		:	dataRd	 = 	 1'b0
;    3182		:	dataRd	 = 	 1'b0
;    3183		:	dataRd	 = 	 1'b0
;    3184		:	dataRd	 = 	 1'b0
;    3185		:	dataRd	 = 	 1'b0
;    3186		:	dataRd	 = 	 1'b0
;    3187		:	dataRd	 = 	 1'b0
;    3188		:	dataRd	 = 	 1'b0
;    3189		:	dataRd	 = 	 1'b0
;    3190		:	dataRd	 = 	 1'b0
;    3191		:	dataRd	 = 	 1'b0
;    3192		:	dataRd	 = 	 1'b0
;    3193		:	dataRd	 = 	 1'b0
;    3194		:	dataRd	 = 	 1'b0
;    3195		:	dataRd	 = 	 1'b0
;    3196		:	dataRd	 = 	 1'b0
;    3197		:	dataRd	 = 	 1'b0
;    3198		:	dataRd	 = 	 1'b0
;    3199		:	dataRd	 = 	 1'b0
;    3200		:	dataRd	 = 	 1'b0
;    3201		:	dataRd	 = 	 1'b0
;    3202		:	dataRd	 = 	 1'b0
;    3203		:	dataRd	 = 	 1'b0
;    3204		:	dataRd	 = 	 1'b0
;    3205		:	dataRd	 = 	 1'b0
;    3206		:	dataRd	 = 	 1'b0
;    3207		:	dataRd	 = 	 1'b0
;    3208		:	dataRd	 = 	 1'b0
;    3209		:	dataRd	 = 	 1'b0
;    3210		:	dataRd	 = 	 1'b0
;    3211		:	dataRd	 = 	 1'b0
;    3212		:	dataRd	 = 	 1'b0
;    3213		:	dataRd	 = 	 1'b0
;    3214		:	dataRd	 = 	 1'b0
;    3215		:	dataRd	 = 	 1'b0
;    3216		:	dataRd	 = 	 1'b0
;    3217		:	dataRd	 = 	 1'b0
;    3218		:	dataRd	 = 	 1'b0
;    3219		:	dataRd	 = 	 1'b0
;    3220		:	dataRd	 = 	 1'b0
;    3221		:	dataRd	 = 	 1'b0
;    3222		:	dataRd	 = 	 1'b0
;    3223		:	dataRd	 = 	 1'b0
;    3224		:	dataRd	 = 	 1'b0
;    3225		:	dataRd	 = 	 1'b0
;    3226		:	dataRd	 = 	 1'b0
;    3227		:	dataRd	 = 	 1'b0
;    3228		:	dataRd	 = 	 1'b0
;    3229		:	dataRd	 = 	 1'b0
;    3230		:	dataRd	 = 	 1'b0
;    3231		:	dataRd	 = 	 1'b0
;    3232		:	dataRd	 = 	 1'b0
;    3233		:	dataRd	 = 	 1'b0
;    3234		:	dataRd	 = 	 1'b0
;    3235		:	dataRd	 = 	 1'b0
;    3236		:	dataRd	 = 	 1'b0
;    3237		:	dataRd	 = 	 1'b0
;    3238		:	dataRd	 = 	 1'b0
;    3239		:	dataRd	 = 	 1'b0
;    3240		:	dataRd	 = 	 1'b0
;    3241		:	dataRd	 = 	 1'b0
;    3242		:	dataRd	 = 	 1'b0
;    3243		:	dataRd	 = 	 1'b0
;    3244		:	dataRd	 = 	 1'b1
;    3245		:	dataRd	 = 	 1'b0
;    3246		:	dataRd	 = 	 1'b0
;    3247		:	dataRd	 = 	 1'b0
;    3248		:	dataRd	 = 	 1'b0
;    3249		:	dataRd	 = 	 1'b0
;    3250		:	dataRd	 = 	 1'b0
;    3251		:	dataRd	 = 	 1'b0
;    3252		:	dataRd	 = 	 1'b0
;    3253		:	dataRd	 = 	 1'b0
;    3254		:	dataRd	 = 	 1'b0
;    3255		:	dataRd	 = 	 1'b0
;    3256		:	dataRd	 = 	 1'b0
;    3257		:	dataRd	 = 	 1'b0
;    3258		:	dataRd	 = 	 1'b0
;    3259		:	dataRd	 = 	 1'b0
;    3260		:	dataRd	 = 	 1'b0
;    3261		:	dataRd	 = 	 1'b0
;    3262		:	dataRd	 = 	 1'b0
;    3263		:	dataRd	 = 	 1'b0
;    3264		:	dataRd	 = 	 1'b0
;    3265		:	dataRd	 = 	 1'b0
;    3266		:	dataRd	 = 	 1'b0
;    3267		:	dataRd	 = 	 1'b0
;    3268		:	dataRd	 = 	 1'b0
;    3269		:	dataRd	 = 	 1'b0
;    3270		:	dataRd	 = 	 1'b0
;    3271		:	dataRd	 = 	 1'b0
;    3272		:	dataRd	 = 	 1'b0
;    3273		:	dataRd	 = 	 1'b0
;    3274		:	dataRd	 = 	 1'b0
;    3275		:	dataRd	 = 	 1'b0
;    3276		:	dataRd	 = 	 1'b0
;    3277		:	dataRd	 = 	 1'b0
;    3278		:	dataRd	 = 	 1'b0
;    3279		:	dataRd	 = 	 1'b0
;    3280		:	dataRd	 = 	 1'b0
;    3281		:	dataRd	 = 	 1'b0
;    3282		:	dataRd	 = 	 1'b0
;    3283		:	dataRd	 = 	 1'b0
;    3284		:	dataRd	 = 	 1'b0
;    3285		:	dataRd	 = 	 1'b0
;    3286		:	dataRd	 = 	 1'b0
;    3287		:	dataRd	 = 	 1'b0
;    3288		:	dataRd	 = 	 1'b0
;    3289		:	dataRd	 = 	 1'b0
;    3290		:	dataRd	 = 	 1'b0
;    3291		:	dataRd	 = 	 1'b0
;    3292		:	dataRd	 = 	 1'b0
;    3293		:	dataRd	 = 	 1'b0
;    3294		:	dataRd	 = 	 1'b0
;    3295		:	dataRd	 = 	 1'b0
;    3296		:	dataRd	 = 	 1'b0
;    3297		:	dataRd	 = 	 1'b0
;    3298		:	dataRd	 = 	 1'b0
;    3299		:	dataRd	 = 	 1'b0
;    3300		:	dataRd	 = 	 1'b0
;    3301		:	dataRd	 = 	 1'b0
;    3302		:	dataRd	 = 	 1'b0
;    3303		:	dataRd	 = 	 1'b0
;    3304		:	dataRd	 = 	 1'b0
;    3305		:	dataRd	 = 	 1'b0
;    3306		:	dataRd	 = 	 1'b0
;    3307		:	dataRd	 = 	 1'b0
;    3308		:	dataRd	 = 	 1'b0
;    3309		:	dataRd	 = 	 1'b0
;    3310		:	dataRd	 = 	 1'b0
;    3311		:	dataRd	 = 	 1'b1
;    3312		:	dataRd	 = 	 1'b0
;    3313		:	dataRd	 = 	 1'b0
;    3314		:	dataRd	 = 	 1'b0
;    3315		:	dataRd	 = 	 1'b0
;    3316		:	dataRd	 = 	 1'b0
;    3317		:	dataRd	 = 	 1'b0
;    3318		:	dataRd	 = 	 1'b0
;    3319		:	dataRd	 = 	 1'b0
;    3320		:	dataRd	 = 	 1'b0
;    3321		:	dataRd	 = 	 1'b0
;    3322		:	dataRd	 = 	 1'b0
;    3323		:	dataRd	 = 	 1'b0
;    3324		:	dataRd	 = 	 1'b0
;    3325		:	dataRd	 = 	 1'b0
;    3326		:	dataRd	 = 	 1'b0
;    3327		:	dataRd	 = 	 1'b0
;    3328		:	dataRd	 = 	 1'b0
;    3329		:	dataRd	 = 	 1'b0
;    3330		:	dataRd	 = 	 1'b0
;    3331		:	dataRd	 = 	 1'b0
;    3332		:	dataRd	 = 	 1'b0
;    3333		:	dataRd	 = 	 1'b0
;    3334		:	dataRd	 = 	 1'b0
;    3335		:	dataRd	 = 	 1'b0
;    3336		:	dataRd	 = 	 1'b0
;    3337		:	dataRd	 = 	 1'b0
;    3338		:	dataRd	 = 	 1'b0
;    3339		:	dataRd	 = 	 1'b0
;    3340		:	dataRd	 = 	 1'b0
;    3341		:	dataRd	 = 	 1'b0
;    3342		:	dataRd	 = 	 1'b0
;    3343		:	dataRd	 = 	 1'b0
;    3344		:	dataRd	 = 	 1'b0
;    3345		:	dataRd	 = 	 1'b0
;    3346		:	dataRd	 = 	 1'b0
;    3347		:	dataRd	 = 	 1'b0
;    3348		:	dataRd	 = 	 1'b0
;    3349		:	dataRd	 = 	 1'b0
;    3350		:	dataRd	 = 	 1'b0
;    3351		:	dataRd	 = 	 1'b0
;    3352		:	dataRd	 = 	 1'b0
;    3353		:	dataRd	 = 	 1'b0
;    3354		:	dataRd	 = 	 1'b0
;    3355		:	dataRd	 = 	 1'b0
;    3356		:	dataRd	 = 	 1'b0
;    3357		:	dataRd	 = 	 1'b0
;    3358		:	dataRd	 = 	 1'b0
;    3359		:	dataRd	 = 	 1'b0
;    3360		:	dataRd	 = 	 1'b0
;    3361		:	dataRd	 = 	 1'b0
;    3362		:	dataRd	 = 	 1'b0
;    3363		:	dataRd	 = 	 1'b0
;    3364		:	dataRd	 = 	 1'b0
;    3365		:	dataRd	 = 	 1'b0
;    3366		:	dataRd	 = 	 1'b0
;    3367		:	dataRd	 = 	 1'b0
;    3368		:	dataRd	 = 	 1'b0
;    3369		:	dataRd	 = 	 1'b0
;    3370		:	dataRd	 = 	 1'b0
;    3371		:	dataRd	 = 	 1'b0
;    3372		:	dataRd	 = 	 1'b0
;    3373		:	dataRd	 = 	 1'b0
;    3374		:	dataRd	 = 	 1'b0
;    3375		:	dataRd	 = 	 1'b0
;    3376		:	dataRd	 = 	 1'b0
;    3377		:	dataRd	 = 	 1'b0
;    3378		:	dataRd	 = 	 1'b0
;    3379		:	dataRd	 = 	 1'b0
;    3380		:	dataRd	 = 	 1'b0
;    3381		:	dataRd	 = 	 1'b0
;    3382		:	dataRd	 = 	 1'b0
;    3383		:	dataRd	 = 	 1'b0
;    3384		:	dataRd	 = 	 1'b0
;    3385		:	dataRd	 = 	 1'b0
;    3386		:	dataRd	 = 	 1'b0
;    3387		:	dataRd	 = 	 1'b0
;    3388		:	dataRd	 = 	 1'b0
;    3389		:	dataRd	 = 	 1'b0
;    3390		:	dataRd	 = 	 1'b0
;    3391		:	dataRd	 = 	 1'b0
;    3392		:	dataRd	 = 	 1'b0
;    3393		:	dataRd	 = 	 1'b0
;    3394		:	dataRd	 = 	 1'b0
;    3395		:	dataRd	 = 	 1'b0
;    3396		:	dataRd	 = 	 1'b0
;    3397		:	dataRd	 = 	 1'b0
;    3398		:	dataRd	 = 	 1'b0
;    3399		:	dataRd	 = 	 1'b0
;    3400		:	dataRd	 = 	 1'b0
;    3401		:	dataRd	 = 	 1'b0
;    3402		:	dataRd	 = 	 1'b0
;    3403		:	dataRd	 = 	 1'b0
;    3404		:	dataRd	 = 	 1'b0
;    3405		:	dataRd	 = 	 1'b0
;    3406		:	dataRd	 = 	 1'b0
;    3407		:	dataRd	 = 	 1'b0
;    3408		:	dataRd	 = 	 1'b0
;    3409		:	dataRd	 = 	 1'b0
;    3410		:	dataRd	 = 	 1'b0
;    3411		:	dataRd	 = 	 1'b0
;    3412		:	dataRd	 = 	 1'b0
;    3413		:	dataRd	 = 	 1'b0
;    3414		:	dataRd	 = 	 1'b0
;    3415		:	dataRd	 = 	 1'b0
;    3416		:	dataRd	 = 	 1'b0
;    3417		:	dataRd	 = 	 1'b0
;    3418		:	dataRd	 = 	 1'b0
;    3419		:	dataRd	 = 	 1'b0
;    3420		:	dataRd	 = 	 1'b0
;    3421		:	dataRd	 = 	 1'b0
;    3422		:	dataRd	 = 	 1'b0
;    3423		:	dataRd	 = 	 1'b0
;    3424		:	dataRd	 = 	 1'b0
;    3425		:	dataRd	 = 	 1'b0
;    3426		:	dataRd	 = 	 1'b0
;    3427		:	dataRd	 = 	 1'b0
;    3428		:	dataRd	 = 	 1'b0
;    3429		:	dataRd	 = 	 1'b0
;    3430		:	dataRd	 = 	 1'b0
;    3431		:	dataRd	 = 	 1'b0
;    3432		:	dataRd	 = 	 1'b0
;    3433		:	dataRd	 = 	 1'b0
;    3434		:	dataRd	 = 	 1'b0
;    3435		:	dataRd	 = 	 1'b0
;    3436		:	dataRd	 = 	 1'b0
;    3437		:	dataRd	 = 	 1'b0
;    3438		:	dataRd	 = 	 1'b0
;    3439		:	dataRd	 = 	 1'b0
;    3440		:	dataRd	 = 	 1'b0
;    3441		:	dataRd	 = 	 1'b0
;    3442		:	dataRd	 = 	 1'b0
;    3443		:	dataRd	 = 	 1'b0
;    3444		:	dataRd	 = 	 1'b1
;    3445		:	dataRd	 = 	 1'b0
;    3446		:	dataRd	 = 	 1'b0
;    3447		:	dataRd	 = 	 1'b0
;    3448		:	dataRd	 = 	 1'b0
;    3449		:	dataRd	 = 	 1'b0
;    3450		:	dataRd	 = 	 1'b0
;    3451		:	dataRd	 = 	 1'b0
;    3452		:	dataRd	 = 	 1'b1
;    3453		:	dataRd	 = 	 1'b0
;    3454		:	dataRd	 = 	 1'b0
;    3455		:	dataRd	 = 	 1'b0
;    3456		:	dataRd	 = 	 1'b0
;    3457		:	dataRd	 = 	 1'b0
;    3458		:	dataRd	 = 	 1'b0
;    3459		:	dataRd	 = 	 1'b0
;    3460		:	dataRd	 = 	 1'b1
;    3461		:	dataRd	 = 	 1'b0
;    3462		:	dataRd	 = 	 1'b0
;    3463		:	dataRd	 = 	 1'b0
;    3464		:	dataRd	 = 	 1'b0
;    3465		:	dataRd	 = 	 1'b0
;    3466		:	dataRd	 = 	 1'b0
;    3467		:	dataRd	 = 	 1'b0
;    3468		:	dataRd	 = 	 1'b1
;    3469		:	dataRd	 = 	 1'b0
;    3470		:	dataRd	 = 	 1'b0
;    3471		:	dataRd	 = 	 1'b1
;    3472		:	dataRd	 = 	 1'b0
;    3473		:	dataRd	 = 	 1'b0
;    3474		:	dataRd	 = 	 1'b1
;    3475		:	dataRd	 = 	 1'b0
;    3476		:	dataRd	 = 	 1'b0
;    3477		:	dataRd	 = 	 1'b0
;    3478		:	dataRd	 = 	 1'b0
;    3479		:	dataRd	 = 	 1'b0
;    3480		:	dataRd	 = 	 1'b0
;    3481		:	dataRd	 = 	 1'b0
;    3482		:	dataRd	 = 	 1'b0
;    3483		:	dataRd	 = 	 1'b0
;    3484		:	dataRd	 = 	 1'b0
;    3485		:	dataRd	 = 	 1'b0
;    3486		:	dataRd	 = 	 1'b0
;    3487		:	dataRd	 = 	 1'b0
;    3488		:	dataRd	 = 	 1'b1
;    3489		:	dataRd	 = 	 1'b0
;    3490		:	dataRd	 = 	 1'b0
;    3491		:	dataRd	 = 	 1'b0
;    3492		:	dataRd	 = 	 1'b0
;    3493		:	dataRd	 = 	 1'b0
;    3494		:	dataRd	 = 	 1'b0
;    3495		:	dataRd	 = 	 1'b1
;    3496		:	dataRd	 = 	 1'b0
;    3497		:	dataRd	 = 	 1'b0
;    3498		:	dataRd	 = 	 1'b1
;    3499		:	dataRd	 = 	 1'b0
;    3500		:	dataRd	 = 	 1'b0
;    3501		:	dataRd	 = 	 1'b0
;    3502		:	dataRd	 = 	 1'b0
;    3503		:	dataRd	 = 	 1'b0
;    3504		:	dataRd	 = 	 1'b0
;    3505		:	dataRd	 = 	 1'b0
;    3506		:	dataRd	 = 	 1'b0
;    3507		:	dataRd	 = 	 1'b0
;    3508		:	dataRd	 = 	 1'b0
;    3509		:	dataRd	 = 	 1'b0
;    3510		:	dataRd	 = 	 1'b0
;    3511		:	dataRd	 = 	 1'b0
;    3512		:	dataRd	 = 	 1'b0
;    3513		:	dataRd	 = 	 1'b0
;    3514		:	dataRd	 = 	 1'b0
;    3515		:	dataRd	 = 	 1'b0
;    3516		:	dataRd	 = 	 1'b0
;    3517		:	dataRd	 = 	 1'b0
;    3518		:	dataRd	 = 	 1'b0
;    3519		:	dataRd	 = 	 1'b1
;    3520		:	dataRd	 = 	 1'b0
;    3521		:	dataRd	 = 	 1'b0
;    3522		:	dataRd	 = 	 1'b0
;    3523		:	dataRd	 = 	 1'b0
;    3524		:	dataRd	 = 	 1'b0
;    3525		:	dataRd	 = 	 1'b0
;    3526		:	dataRd	 = 	 1'b0
;    3527		:	dataRd	 = 	 1'b1
;    3528		:	dataRd	 = 	 1'b0
;    3529		:	dataRd	 = 	 1'b0
;    3530		:	dataRd	 = 	 1'b1
;    3531		:	dataRd	 = 	 1'b0
;    3532		:	dataRd	 = 	 1'b0
;    3533		:	dataRd	 = 	 1'b0
;    3534		:	dataRd	 = 	 1'b0
;    3535		:	dataRd	 = 	 1'b0
;    3536		:	dataRd	 = 	 1'b0
;    3537		:	dataRd	 = 	 1'b0
;    3538		:	dataRd	 = 	 1'b0
;    3539		:	dataRd	 = 	 1'b0
;    3540		:	dataRd	 = 	 1'b0
;    3541		:	dataRd	 = 	 1'b0
;    3542		:	dataRd	 = 	 1'b0
;    3543		:	dataRd	 = 	 1'b0
;    3544		:	dataRd	 = 	 1'b0
;    3545		:	dataRd	 = 	 1'b0
;    3546		:	dataRd	 = 	 1'b1
;    3547		:	dataRd	 = 	 1'b0
;    3548		:	dataRd	 = 	 1'b0
;    3549		:	dataRd	 = 	 1'b0
;    3550		:	dataRd	 = 	 1'b0
;    3551		:	dataRd	 = 	 1'b0
;    3552		:	dataRd	 = 	 1'b0
;    3553		:	dataRd	 = 	 1'b0
;    3554		:	dataRd	 = 	 1'b0
;    3555		:	dataRd	 = 	 1'b0
;    3556		:	dataRd	 = 	 1'b0
;    3557		:	dataRd	 = 	 1'b0
;    3558		:	dataRd	 = 	 1'b0
;    3559		:	dataRd	 = 	 1'b0
;    3560		:	dataRd	 = 	 1'b0
;    3561		:	dataRd	 = 	 1'b0
;    3562		:	dataRd	 = 	 1'b1
;    3563		:	dataRd	 = 	 1'b0
;    3564		:	dataRd	 = 	 1'b0
;    3565		:	dataRd	 = 	 1'b0
;    3566		:	dataRd	 = 	 1'b0
;    3567		:	dataRd	 = 	 1'b0
;    3568		:	dataRd	 = 	 1'b0
;    3569		:	dataRd	 = 	 1'b0
;    3570		:	dataRd	 = 	 1'b0
;    3571		:	dataRd	 = 	 1'b0
;    3572		:	dataRd	 = 	 1'b0
;    3573		:	dataRd	 = 	 1'b0
;    3574		:	dataRd	 = 	 1'b0
;    3575		:	dataRd	 = 	 1'b0
;    3576		:	dataRd	 = 	 1'b0
;    3577		:	dataRd	 = 	 1'b0
;    3578		:	dataRd	 = 	 1'b1
;    3579		:	dataRd	 = 	 1'b0
;    3580		:	dataRd	 = 	 1'b0
;    3581		:	dataRd	 = 	 1'b0
;    3582		:	dataRd	 = 	 1'b0
;    3583		:	dataRd	 = 	 1'b0
;    3584		:	dataRd	 = 	 1'b0
;    3585		:	dataRd	 = 	 1'b0
;    3586		:	dataRd	 = 	 1'b0
;    3587		:	dataRd	 = 	 1'b0
;    3588		:	dataRd	 = 	 1'b0
;    3589		:	dataRd	 = 	 1'b0
;    3590		:	dataRd	 = 	 1'b0
;    3591		:	dataRd	 = 	 1'b0
;    3592		:	dataRd	 = 	 1'b0
;    3593		:	dataRd	 = 	 1'b0
;    3594		:	dataRd	 = 	 1'b1
;    3595		:	dataRd	 = 	 1'b0
;    3596		:	dataRd	 = 	 1'b0
;    3597		:	dataRd	 = 	 1'b0
;    3598		:	dataRd	 = 	 1'b0
;    3599		:	dataRd	 = 	 1'b0
;    3600		:	dataRd	 = 	 1'b0
;    3601		:	dataRd	 = 	 1'b0
;    3602		:	dataRd	 = 	 1'b0
;    3603		:	dataRd	 = 	 1'b0
;    3604		:	dataRd	 = 	 1'b0
;    3605		:	dataRd	 = 	 1'b0
;    3606		:	dataRd	 = 	 1'b0
;    3607		:	dataRd	 = 	 1'b0
;    3608		:	dataRd	 = 	 1'b0
;    3609		:	dataRd	 = 	 1'b0
;    3610		:	dataRd	 = 	 1'b1
;    3611		:	dataRd	 = 	 1'b0
;    3612		:	dataRd	 = 	 1'b0
;    3613		:	dataRd	 = 	 1'b0
;    3614		:	dataRd	 = 	 1'b0
;    3615		:	dataRd	 = 	 1'b0
;    3616		:	dataRd	 = 	 1'b0
;    3617		:	dataRd	 = 	 1'b0
;    3618		:	dataRd	 = 	 1'b0
;    3619		:	dataRd	 = 	 1'b0
;    3620		:	dataRd	 = 	 1'b0
;    3621		:	dataRd	 = 	 1'b0
;    3622		:	dataRd	 = 	 1'b0
;    3623		:	dataRd	 = 	 1'b0
;    3624		:	dataRd	 = 	 1'b0
;    3625		:	dataRd	 = 	 1'b0
;    3626		:	dataRd	 = 	 1'b1
;    3627		:	dataRd	 = 	 1'b0
;    3628		:	dataRd	 = 	 1'b0
;    3629		:	dataRd	 = 	 1'b0
;    3630		:	dataRd	 = 	 1'b0
;    3631		:	dataRd	 = 	 1'b0
;    3632		:	dataRd	 = 	 1'b0
;    3633		:	dataRd	 = 	 1'b0
;    3634		:	dataRd	 = 	 1'b0
;    3635		:	dataRd	 = 	 1'b0
;    3636		:	dataRd	 = 	 1'b0
;    3637		:	dataRd	 = 	 1'b0
;    3638		:	dataRd	 = 	 1'b0
;    3639		:	dataRd	 = 	 1'b0
;    3640		:	dataRd	 = 	 1'b0
;    3641		:	dataRd	 = 	 1'b0
;    3642		:	dataRd	 = 	 1'b1
;    3643		:	dataRd	 = 	 1'b0
;    3644		:	dataRd	 = 	 1'b0
;    3645		:	dataRd	 = 	 1'b0
;    3646		:	dataRd	 = 	 1'b0
;    3647		:	dataRd	 = 	 1'b0
;    3648		:	dataRd	 = 	 1'b0
;    3649		:	dataRd	 = 	 1'b0
;    3650		:	dataRd	 = 	 1'b0
;    3651		:	dataRd	 = 	 1'b0
;    3652		:	dataRd	 = 	 1'b0
;    3653		:	dataRd	 = 	 1'b0
;    3654		:	dataRd	 = 	 1'b0
;    3655		:	dataRd	 = 	 1'b0
;    3656		:	dataRd	 = 	 1'b0
;    3657		:	dataRd	 = 	 1'b0
;    3658		:	dataRd	 = 	 1'b1
;    3659		:	dataRd	 = 	 1'b0
;    3660		:	dataRd	 = 	 1'b0
;    3661		:	dataRd	 = 	 1'b0
;    3662		:	dataRd	 = 	 1'b0
;    3663		:	dataRd	 = 	 1'b0
;    3664		:	dataRd	 = 	 1'b0
;    3665		:	dataRd	 = 	 1'b0
;    3666		:	dataRd	 = 	 1'b0
;    3667		:	dataRd	 = 	 1'b0
;    3668		:	dataRd	 = 	 1'b0
;    3669		:	dataRd	 = 	 1'b0
;    3670		:	dataRd	 = 	 1'b0
;    3671		:	dataRd	 = 	 1'b0
;    3672		:	dataRd	 = 	 1'b0
;    3673		:	dataRd	 = 	 1'b0
;    3674		:	dataRd	 = 	 1'b1
;    3675		:	dataRd	 = 	 1'b0
;    3676		:	dataRd	 = 	 1'b0
;    3677		:	dataRd	 = 	 1'b0
;    3678		:	dataRd	 = 	 1'b0
;    3679		:	dataRd	 = 	 1'b0
;    3680		:	dataRd	 = 	 1'b0
;    3681		:	dataRd	 = 	 1'b0
;    3682		:	dataRd	 = 	 1'b0
;    3683		:	dataRd	 = 	 1'b0
;    3684		:	dataRd	 = 	 1'b0
;    3685		:	dataRd	 = 	 1'b0
;    3686		:	dataRd	 = 	 1'b0
;    3687		:	dataRd	 = 	 1'b0
;    3688		:	dataRd	 = 	 1'b0
;    3689		:	dataRd	 = 	 1'b0
;    3690		:	dataRd	 = 	 1'b1
;    3691		:	dataRd	 = 	 1'b0
;    3692		:	dataRd	 = 	 1'b0
;    3693		:	dataRd	 = 	 1'b0
;    3694		:	dataRd	 = 	 1'b0
;    3695		:	dataRd	 = 	 1'b0
;    3696		:	dataRd	 = 	 1'b0
;    3697		:	dataRd	 = 	 1'b0
;    3698		:	dataRd	 = 	 1'b0
;    3699		:	dataRd	 = 	 1'b0
;    3700		:	dataRd	 = 	 1'b0
;    3701		:	dataRd	 = 	 1'b0
;    3702		:	dataRd	 = 	 1'b0
;    3703		:	dataRd	 = 	 1'b0
;    3704		:	dataRd	 = 	 1'b0
;    3705		:	dataRd	 = 	 1'b0
;    3706		:	dataRd	 = 	 1'b1
;    3707		:	dataRd	 = 	 1'b0
;    3708		:	dataRd	 = 	 1'b0
;    3709		:	dataRd	 = 	 1'b0
;    3710		:	dataRd	 = 	 1'b0
;    3711		:	dataRd	 = 	 1'b0
;    3712		:	dataRd	 = 	 1'b0
;    3713		:	dataRd	 = 	 1'b0
;    3714		:	dataRd	 = 	 1'b0
;    3715		:	dataRd	 = 	 1'b0
;    3716		:	dataRd	 = 	 1'b0
;    3717		:	dataRd	 = 	 1'b0
;    3718		:	dataRd	 = 	 1'b0
;    3719		:	dataRd	 = 	 1'b0
;    3720		:	dataRd	 = 	 1'b0
;    3721		:	dataRd	 = 	 1'b0
;    3722		:	dataRd	 = 	 1'b1
;    3723		:	dataRd	 = 	 1'b0
;    3724		:	dataRd	 = 	 1'b0
;    3725		:	dataRd	 = 	 1'b0
;    3726		:	dataRd	 = 	 1'b0
;    3727		:	dataRd	 = 	 1'b0
;    3728		:	dataRd	 = 	 1'b0
;    3729		:	dataRd	 = 	 1'b0
;    3730		:	dataRd	 = 	 1'b0
;    3731		:	dataRd	 = 	 1'b0
;    3732		:	dataRd	 = 	 1'b0
;    3733		:	dataRd	 = 	 1'b0
;    3734		:	dataRd	 = 	 1'b0
;    3735		:	dataRd	 = 	 1'b0
;    3736		:	dataRd	 = 	 1'b0
;    3737		:	dataRd	 = 	 1'b0
;    3738		:	dataRd	 = 	 1'b1
;    3739		:	dataRd	 = 	 1'b0
;    3740		:	dataRd	 = 	 1'b0
;    3741		:	dataRd	 = 	 1'b0
;    3742		:	dataRd	 = 	 1'b0
;    3743		:	dataRd	 = 	 1'b0
;    3744		:	dataRd	 = 	 1'b0
;    3745		:	dataRd	 = 	 1'b0
;    3746		:	dataRd	 = 	 1'b0
;    3747		:	dataRd	 = 	 1'b0
;    3748		:	dataRd	 = 	 1'b0
;    3749		:	dataRd	 = 	 1'b0
;    3750		:	dataRd	 = 	 1'b0
;    3751		:	dataRd	 = 	 1'b0
;    3752		:	dataRd	 = 	 1'b0
;    3753		:	dataRd	 = 	 1'b0
;    3754		:	dataRd	 = 	 1'b1
;    3755		:	dataRd	 = 	 1'b0
;    3756		:	dataRd	 = 	 1'b0
;    3757		:	dataRd	 = 	 1'b0
;    3758		:	dataRd	 = 	 1'b0
;    3759		:	dataRd	 = 	 1'b0
;    3760		:	dataRd	 = 	 1'b0
;    3761		:	dataRd	 = 	 1'b0
;    3762		:	dataRd	 = 	 1'b0
;    3763		:	dataRd	 = 	 1'b0
;    3764		:	dataRd	 = 	 1'b0
;    3765		:	dataRd	 = 	 1'b0
;    3766		:	dataRd	 = 	 1'b0
;    3767		:	dataRd	 = 	 1'b0
;    3768		:	dataRd	 = 	 1'b0
;    3769		:	dataRd	 = 	 1'b0
;    3770		:	dataRd	 = 	 1'b1
;    3771		:	dataRd	 = 	 1'b0
;    3772		:	dataRd	 = 	 1'b0
;    3773		:	dataRd	 = 	 1'b0
;    3774		:	dataRd	 = 	 1'b0
;    3775		:	dataRd	 = 	 1'b0
;    3776		:	dataRd	 = 	 1'b0
;    3777		:	dataRd	 = 	 1'b0
;    3778		:	dataRd	 = 	 1'b0
;    3779		:	dataRd	 = 	 1'b0
;    3780		:	dataRd	 = 	 1'b0
;    3781		:	dataRd	 = 	 1'b0
;    3782		:	dataRd	 = 	 1'b0
;    3783		:	dataRd	 = 	 1'b0
;    3784		:	dataRd	 = 	 1'b0
;    3785		:	dataRd	 = 	 1'b0
;    3786		:	dataRd	 = 	 1'b1
;    3787		:	dataRd	 = 	 1'b0
;    3788		:	dataRd	 = 	 1'b0
;    3789		:	dataRd	 = 	 1'b0
;    3790		:	dataRd	 = 	 1'b0
;    3791		:	dataRd	 = 	 1'b0
;    3792		:	dataRd	 = 	 1'b0
;    3793		:	dataRd	 = 	 1'b0
;    3794		:	dataRd	 = 	 1'b0
;    3795		:	dataRd	 = 	 1'b0
;    3796		:	dataRd	 = 	 1'b0
;    3797		:	dataRd	 = 	 1'b0
;    3798		:	dataRd	 = 	 1'b0
;    3799		:	dataRd	 = 	 1'b0
;    3800		:	dataRd	 = 	 1'b0
;    3801		:	dataRd	 = 	 1'b0
;    3802		:	dataRd	 = 	 1'b1
;    3803		:	dataRd	 = 	 1'b0
;    3804		:	dataRd	 = 	 1'b0
;    3805		:	dataRd	 = 	 1'b0
;    3806		:	dataRd	 = 	 1'b0
;    3807		:	dataRd	 = 	 1'b0
;    3808		:	dataRd	 = 	 1'b0
;    3809		:	dataRd	 = 	 1'b0
;    3810		:	dataRd	 = 	 1'b0
;    3811		:	dataRd	 = 	 1'b0
;    3812		:	dataRd	 = 	 1'b0
;    3813		:	dataRd	 = 	 1'b0
;    3814		:	dataRd	 = 	 1'b0
;    3815		:	dataRd	 = 	 1'b0
;    3816		:	dataRd	 = 	 1'b0
;    3817		:	dataRd	 = 	 1'b0
;    3818		:	dataRd	 = 	 1'b1
;    3819		:	dataRd	 = 	 1'b0
;    3820		:	dataRd	 = 	 1'b0
;    3821		:	dataRd	 = 	 1'b0
;    3822		:	dataRd	 = 	 1'b0
;    3823		:	dataRd	 = 	 1'b0
;    3824		:	dataRd	 = 	 1'b0
;    3825		:	dataRd	 = 	 1'b0
;    3826		:	dataRd	 = 	 1'b0
;    3827		:	dataRd	 = 	 1'b0
;    3828		:	dataRd	 = 	 1'b0
;    3829		:	dataRd	 = 	 1'b0
;    3830		:	dataRd	 = 	 1'b0
;    3831		:	dataRd	 = 	 1'b0
;    3832		:	dataRd	 = 	 1'b0
;    3833		:	dataRd	 = 	 1'b0
;    3834		:	dataRd	 = 	 1'b1
;    3835		:	dataRd	 = 	 1'b0
;    3836		:	dataRd	 = 	 1'b0
;    3837		:	dataRd	 = 	 1'b0
;    3838		:	dataRd	 = 	 1'b0
;    3839		:	dataRd	 = 	 1'b0
;    3840		:	dataRd	 = 	 1'b0
;    3841		:	dataRd	 = 	 1'b0
;    3842		:	dataRd	 = 	 1'b0
;    3843		:	dataRd	 = 	 1'b0
;    3844		:	dataRd	 = 	 1'b0
;    3845		:	dataRd	 = 	 1'b0
;    3846		:	dataRd	 = 	 1'b0
;    3847		:	dataRd	 = 	 1'b0
;    3848		:	dataRd	 = 	 1'b0
;    3849		:	dataRd	 = 	 1'b0
;    3850		:	dataRd	 = 	 1'b1
;    3851		:	dataRd	 = 	 1'b0
;    3852		:	dataRd	 = 	 1'b0
;    3853		:	dataRd	 = 	 1'b0
;    3854		:	dataRd	 = 	 1'b0
;    3855		:	dataRd	 = 	 1'b0
;    3856		:	dataRd	 = 	 1'b0
;    3857		:	dataRd	 = 	 1'b0
;    3858		:	dataRd	 = 	 1'b0
;    3859		:	dataRd	 = 	 1'b0
;    3860		:	dataRd	 = 	 1'b0
;    3861		:	dataRd	 = 	 1'b0
;    3862		:	dataRd	 = 	 1'b0
;    3863		:	dataRd	 = 	 1'b0
;    3864		:	dataRd	 = 	 1'b0
;    3865		:	dataRd	 = 	 1'b0
;    3866		:	dataRd	 = 	 1'b1
;    3867		:	dataRd	 = 	 1'b0
;    3868		:	dataRd	 = 	 1'b0
;    3869		:	dataRd	 = 	 1'b0
;    3870		:	dataRd	 = 	 1'b0
;    3871		:	dataRd	 = 	 1'b0
;    3872		:	dataRd	 = 	 1'b0
;    3873		:	dataRd	 = 	 1'b0
;    3874		:	dataRd	 = 	 1'b0
;    3875		:	dataRd	 = 	 1'b0
;    3876		:	dataRd	 = 	 1'b0
;    3877		:	dataRd	 = 	 1'b0
;    3878		:	dataRd	 = 	 1'b0
;    3879		:	dataRd	 = 	 1'b0
;    3880		:	dataRd	 = 	 1'b0
;    3881		:	dataRd	 = 	 1'b0
;    3882		:	dataRd	 = 	 1'b1
;    3883		:	dataRd	 = 	 1'b0
;    3884		:	dataRd	 = 	 1'b0
;    3885		:	dataRd	 = 	 1'b0
;    3886		:	dataRd	 = 	 1'b0
;    3887		:	dataRd	 = 	 1'b0
;    3888		:	dataRd	 = 	 1'b0
;    3889		:	dataRd	 = 	 1'b0
;    3890		:	dataRd	 = 	 1'b0
;    3891		:	dataRd	 = 	 1'b0
;    3892		:	dataRd	 = 	 1'b0
;    3893		:	dataRd	 = 	 1'b0
;    3894		:	dataRd	 = 	 1'b0
;    3895		:	dataRd	 = 	 1'b0
;    3896		:	dataRd	 = 	 1'b0
;    3897		:	dataRd	 = 	 1'b0
;    3898		:	dataRd	 = 	 1'b1
;    3899		:	dataRd	 = 	 1'b0
;    3900		:	dataRd	 = 	 1'b0
;    3901		:	dataRd	 = 	 1'b0
;    3902		:	dataRd	 = 	 1'b0
;    3903		:	dataRd	 = 	 1'b0
;    3904		:	dataRd	 = 	 1'b0
;    3905		:	dataRd	 = 	 1'b0
;    3906		:	dataRd	 = 	 1'b0
;    3907		:	dataRd	 = 	 1'b0
;    3908		:	dataRd	 = 	 1'b0
;    3909		:	dataRd	 = 	 1'b0
;    3910		:	dataRd	 = 	 1'b0
;    3911		:	dataRd	 = 	 1'b0
;    3912		:	dataRd	 = 	 1'b0
;    3913		:	dataRd	 = 	 1'b0
;    3914		:	dataRd	 = 	 1'b1
;    3915		:	dataRd	 = 	 1'b0
;    3916		:	dataRd	 = 	 1'b0
;    3917		:	dataRd	 = 	 1'b0
;    3918		:	dataRd	 = 	 1'b0
;    3919		:	dataRd	 = 	 1'b0
;    3920		:	dataRd	 = 	 1'b0
;    3921		:	dataRd	 = 	 1'b0
;    3922		:	dataRd	 = 	 1'b0
;    3923		:	dataRd	 = 	 1'b0
;    3924		:	dataRd	 = 	 1'b0
;    3925		:	dataRd	 = 	 1'b0
;    3926		:	dataRd	 = 	 1'b0
;    3927		:	dataRd	 = 	 1'b0
;    3928		:	dataRd	 = 	 1'b0
;    3929		:	dataRd	 = 	 1'b0
;    3930		:	dataRd	 = 	 1'b1
;    3931		:	dataRd	 = 	 1'b0
;    3932		:	dataRd	 = 	 1'b0
;    3933		:	dataRd	 = 	 1'b0
;    3934		:	dataRd	 = 	 1'b0
;    3935		:	dataRd	 = 	 1'b0
;    3936		:	dataRd	 = 	 1'b0
;    3937		:	dataRd	 = 	 1'b0
;    3938		:	dataRd	 = 	 1'b0
;    3939		:	dataRd	 = 	 1'b0
;    3940		:	dataRd	 = 	 1'b0
;    3941		:	dataRd	 = 	 1'b0
;    3942		:	dataRd	 = 	 1'b0
;    3943		:	dataRd	 = 	 1'b0
;    3944		:	dataRd	 = 	 1'b0
;    3945		:	dataRd	 = 	 1'b0
;    3946		:	dataRd	 = 	 1'b1
;    3947		:	dataRd	 = 	 1'b0
;    3948		:	dataRd	 = 	 1'b0
;    3949		:	dataRd	 = 	 1'b0
;    3950		:	dataRd	 = 	 1'b0
;    3951		:	dataRd	 = 	 1'b0
;    3952		:	dataRd	 = 	 1'b0
;    3953		:	dataRd	 = 	 1'b0
;    3954		:	dataRd	 = 	 1'b0
;    3955		:	dataRd	 = 	 1'b0
;    3956		:	dataRd	 = 	 1'b0
;    3957		:	dataRd	 = 	 1'b0
;    3958		:	dataRd	 = 	 1'b0
;    3959		:	dataRd	 = 	 1'b0
;    3960		:	dataRd	 = 	 1'b0
;    3961		:	dataRd	 = 	 1'b0
;    3962		:	dataRd	 = 	 1'b1
;    3963		:	dataRd	 = 	 1'b0
;    3964		:	dataRd	 = 	 1'b0
;    3965		:	dataRd	 = 	 1'b0
;    3966		:	dataRd	 = 	 1'b0
;    3967		:	dataRd	 = 	 1'b0
;    3968		:	dataRd	 = 	 1'b0
;    3969		:	dataRd	 = 	 1'b0
;    3970		:	dataRd	 = 	 1'b0
;    3971		:	dataRd	 = 	 1'b0
;    3972		:	dataRd	 = 	 1'b0
;    3973		:	dataRd	 = 	 1'b0
;    3974		:	dataRd	 = 	 1'b0
;    3975		:	dataRd	 = 	 1'b0
;    3976		:	dataRd	 = 	 1'b0
;    3977		:	dataRd	 = 	 1'b0
;    3978		:	dataRd	 = 	 1'b1
;    3979		:	dataRd	 = 	 1'b0
;    3980		:	dataRd	 = 	 1'b0
;    3981		:	dataRd	 = 	 1'b0
;    3982		:	dataRd	 = 	 1'b0
;    3983		:	dataRd	 = 	 1'b0
;    3984		:	dataRd	 = 	 1'b0
;    3985		:	dataRd	 = 	 1'b0
;    3986		:	dataRd	 = 	 1'b0
;    3987		:	dataRd	 = 	 1'b0
;    3988		:	dataRd	 = 	 1'b0
;    3989		:	dataRd	 = 	 1'b0
;    3990		:	dataRd	 = 	 1'b0
;    3991		:	dataRd	 = 	 1'b0
;    3992		:	dataRd	 = 	 1'b0
;    3993		:	dataRd	 = 	 1'b0
;    3994		:	dataRd	 = 	 1'b1
;    3995		:	dataRd	 = 	 1'b0
;    3996		:	dataRd	 = 	 1'b0
;    3997		:	dataRd	 = 	 1'b0
;    3998		:	dataRd	 = 	 1'b0
;    3999		:	dataRd	 = 	 1'b0
;    4000		:	dataRd	 = 	 1'b0
;    4001		:	dataRd	 = 	 1'b0
;    4002		:	dataRd	 = 	 1'b0
;    4003		:	dataRd	 = 	 1'b0
;    4004		:	dataRd	 = 	 1'b0
;    4005		:	dataRd	 = 	 1'b0
;    4006		:	dataRd	 = 	 1'b0
;    4007		:	dataRd	 = 	 1'b0
;    4008		:	dataRd	 = 	 1'b0
;    4009		:	dataRd	 = 	 1'b0
;    4010		:	dataRd	 = 	 1'b1
;    4011		:	dataRd	 = 	 1'b0
;    4012		:	dataRd	 = 	 1'b0
;    4013		:	dataRd	 = 	 1'b0
;    4014		:	dataRd	 = 	 1'b0
;    4015		:	dataRd	 = 	 1'b0
;    4016		:	dataRd	 = 	 1'b0
;    4017		:	dataRd	 = 	 1'b0
;    4018		:	dataRd	 = 	 1'b0
;    4019		:	dataRd	 = 	 1'b0
;    4020		:	dataRd	 = 	 1'b0
;    4021		:	dataRd	 = 	 1'b0
;    4022		:	dataRd	 = 	 1'b0
;    4023		:	dataRd	 = 	 1'b0
;    4024		:	dataRd	 = 	 1'b0
;    4025		:	dataRd	 = 	 1'b0
;    4026		:	dataRd	 = 	 1'b1
;    4027		:	dataRd	 = 	 1'b0
;    4028		:	dataRd	 = 	 1'b0
;    4029		:	dataRd	 = 	 1'b0
;    4030		:	dataRd	 = 	 1'b0
;    4031		:	dataRd	 = 	 1'b0
;    4032		:	dataRd	 = 	 1'b0
;    4033		:	dataRd	 = 	 1'b0
;    4034		:	dataRd	 = 	 1'b0
;    4035		:	dataRd	 = 	 1'b0
;    4036		:	dataRd	 = 	 1'b0
;    4037		:	dataRd	 = 	 1'b0
;    4038		:	dataRd	 = 	 1'b0
;    4039		:	dataRd	 = 	 1'b0
;    4040		:	dataRd	 = 	 1'b0
;    4041		:	dataRd	 = 	 1'b0
;    4042		:	dataRd	 = 	 1'b1
;    4043		:	dataRd	 = 	 1'b0
;    4044		:	dataRd	 = 	 1'b0
;    4045		:	dataRd	 = 	 1'b0
;    4046		:	dataRd	 = 	 1'b0
;    4047		:	dataRd	 = 	 1'b0
;    4048		:	dataRd	 = 	 1'b0
;    4049		:	dataRd	 = 	 1'b0
;    4050		:	dataRd	 = 	 1'b0
;    4051		:	dataRd	 = 	 1'b0
;    4052		:	dataRd	 = 	 1'b0
;    4053		:	dataRd	 = 	 1'b0
;    4054		:	dataRd	 = 	 1'b0
;    4055		:	dataRd	 = 	 1'b0
;    4056		:	dataRd	 = 	 1'b0
;    4057		:	dataRd	 = 	 1'b0
;    4058		:	dataRd	 = 	 1'b1
;    4059		:	dataRd	 = 	 1'b0
;    4060		:	dataRd	 = 	 1'b0
;    4061		:	dataRd	 = 	 1'b0
;    4062		:	dataRd	 = 	 1'b0
;    4063		:	dataRd	 = 	 1'b0
;    4064		:	dataRd	 = 	 1'b0
;    4065		:	dataRd	 = 	 1'b0
;    4066		:	dataRd	 = 	 1'b0
;    4067		:	dataRd	 = 	 1'b0
;    4068		:	dataRd	 = 	 1'b0
;    4069		:	dataRd	 = 	 1'b0
;    4070		:	dataRd	 = 	 1'b0
;    4071		:	dataRd	 = 	 1'b0
;    4072		:	dataRd	 = 	 1'b0
;    4073		:	dataRd	 = 	 1'b0
;    4074		:	dataRd	 = 	 1'b1
;    4075		:	dataRd	 = 	 1'b0
;    4076		:	dataRd	 = 	 1'b0
;    4077		:	dataRd	 = 	 1'b0
;    4078		:	dataRd	 = 	 1'b0
;    4079		:	dataRd	 = 	 1'b0
;    4080		:	dataRd	 = 	 1'b0
;    4081		:	dataRd	 = 	 1'b0
;    4082		:	dataRd	 = 	 1'b0
;    4083		:	dataRd	 = 	 1'b0
;    4084		:	dataRd	 = 	 1'b0
;    4085		:	dataRd	 = 	 1'b0
;    4086		:	dataRd	 = 	 1'b0
;    4087		:	dataRd	 = 	 1'b0
;    4088		:	dataRd	 = 	 1'b0
;    4089		:	dataRd	 = 	 1'b0
;    4090		:	dataRd	 = 	 1'b1
;    4091		:	dataRd	 = 	 1'b0
;    4092		:	dataRd	 = 	 1'b0
;    4093		:	dataRd	 = 	 1'b0
;    4094		:	dataRd	 = 	 1'b0
;    4095		:	dataRd	 = 	 1'b0
;    4096		:	dataRd	 = 	 1'b0
;    4097		:	dataRd	 = 	 1'b0
;    4098		:	dataRd	 = 	 1'b0
;    4099		:	dataRd	 = 	 1'b0
;    4100		:	dataRd	 = 	 1'b0
;    4101		:	dataRd	 = 	 1'b0
;    4102		:	dataRd	 = 	 1'b0
;    4103		:	dataRd	 = 	 1'b0
;    4104		:	dataRd	 = 	 1'b0
;    4105		:	dataRd	 = 	 1'b0
;    4106		:	dataRd	 = 	 1'b1
;    4107		:	dataRd	 = 	 1'b0
;    4108		:	dataRd	 = 	 1'b0
;    4109		:	dataRd	 = 	 1'b0
;    4110		:	dataRd	 = 	 1'b0
;    4111		:	dataRd	 = 	 1'b0
;    4112		:	dataRd	 = 	 1'b0
;    4113		:	dataRd	 = 	 1'b0
;    4114		:	dataRd	 = 	 1'b0
;    4115		:	dataRd	 = 	 1'b0
;    4116		:	dataRd	 = 	 1'b0
;    4117		:	dataRd	 = 	 1'b0
;    4118		:	dataRd	 = 	 1'b0
;    4119		:	dataRd	 = 	 1'b0
;    4120		:	dataRd	 = 	 1'b0
;    4121		:	dataRd	 = 	 1'b0
;    4122		:	dataRd	 = 	 1'b1
;    4123		:	dataRd	 = 	 1'b0
;    4124		:	dataRd	 = 	 1'b0
;    4125		:	dataRd	 = 	 1'b0
;    4126		:	dataRd	 = 	 1'b0
;    4127		:	dataRd	 = 	 1'b0
;    4128		:	dataRd	 = 	 1'b0
;    4129		:	dataRd	 = 	 1'b0
;    4130		:	dataRd	 = 	 1'b0
;    4131		:	dataRd	 = 	 1'b0
;    4132		:	dataRd	 = 	 1'b0
;    4133		:	dataRd	 = 	 1'b0
;    4134		:	dataRd	 = 	 1'b0
;    4135		:	dataRd	 = 	 1'b0
;    4136		:	dataRd	 = 	 1'b0
;    4137		:	dataRd	 = 	 1'b0
;    4138		:	dataRd	 = 	 1'b1
;    4139		:	dataRd	 = 	 1'b0
;    4140		:	dataRd	 = 	 1'b0
;    4141		:	dataRd	 = 	 1'b0
;    4142		:	dataRd	 = 	 1'b0
;    4143		:	dataRd	 = 	 1'b0
;    4144		:	dataRd	 = 	 1'b0
;    4145		:	dataRd	 = 	 1'b0
;    4146		:	dataRd	 = 	 1'b0
;    4147		:	dataRd	 = 	 1'b0
;    4148		:	dataRd	 = 	 1'b0
;    4149		:	dataRd	 = 	 1'b0
;    4150		:	dataRd	 = 	 1'b0
;    4151		:	dataRd	 = 	 1'b0
;    4152		:	dataRd	 = 	 1'b0
;    4153		:	dataRd	 = 	 1'b0
;    4154		:	dataRd	 = 	 1'b1
;    4155		:	dataRd	 = 	 1'b0
;    4156		:	dataRd	 = 	 1'b0
;    4157		:	dataRd	 = 	 1'b0
;    4158		:	dataRd	 = 	 1'b0
;    4159		:	dataRd	 = 	 1'b0
;    4160		:	dataRd	 = 	 1'b0
;    4161		:	dataRd	 = 	 1'b0
;    4162		:	dataRd	 = 	 1'b0
;    4163		:	dataRd	 = 	 1'b0
;    4164		:	dataRd	 = 	 1'b0
;    4165		:	dataRd	 = 	 1'b0
;    4166		:	dataRd	 = 	 1'b0
;    4167		:	dataRd	 = 	 1'b0
;    4168		:	dataRd	 = 	 1'b0
;    4169		:	dataRd	 = 	 1'b0
;    4170		:	dataRd	 = 	 1'b1
;    4171		:	dataRd	 = 	 1'b0
;    4172		:	dataRd	 = 	 1'b0
;    4173		:	dataRd	 = 	 1'b0
;    4174		:	dataRd	 = 	 1'b0
;    4175		:	dataRd	 = 	 1'b0
;    4176		:	dataRd	 = 	 1'b0
;    4177		:	dataRd	 = 	 1'b0
;    4178		:	dataRd	 = 	 1'b0
;    4179		:	dataRd	 = 	 1'b0
;    4180		:	dataRd	 = 	 1'b0
;    4181		:	dataRd	 = 	 1'b0
;    4182		:	dataRd	 = 	 1'b0
;    4183		:	dataRd	 = 	 1'b0
;    4184		:	dataRd	 = 	 1'b0
;    4185		:	dataRd	 = 	 1'b0
;    4186		:	dataRd	 = 	 1'b1
;    4187		:	dataRd	 = 	 1'b0
;    4188		:	dataRd	 = 	 1'b0
;    4189		:	dataRd	 = 	 1'b0
;    4190		:	dataRd	 = 	 1'b0
;    4191		:	dataRd	 = 	 1'b0
;    4192		:	dataRd	 = 	 1'b0
;    4193		:	dataRd	 = 	 1'b0
;    4194		:	dataRd	 = 	 1'b0
;    4195		:	dataRd	 = 	 1'b0
;    4196		:	dataRd	 = 	 1'b0
;    4197		:	dataRd	 = 	 1'b0
;    4198		:	dataRd	 = 	 1'b0
;    4199		:	dataRd	 = 	 1'b0
;    4200		:	dataRd	 = 	 1'b0
;    4201		:	dataRd	 = 	 1'b0
;    4202		:	dataRd	 = 	 1'b1
;    4203		:	dataRd	 = 	 1'b0
;    4204		:	dataRd	 = 	 1'b0
;    4205		:	dataRd	 = 	 1'b0
;    4206		:	dataRd	 = 	 1'b0
;    4207		:	dataRd	 = 	 1'b0
;    4208		:	dataRd	 = 	 1'b0
;    4209		:	dataRd	 = 	 1'b0
;    4210		:	dataRd	 = 	 1'b0
;    4211		:	dataRd	 = 	 1'b0
;    4212		:	dataRd	 = 	 1'b0
;    4213		:	dataRd	 = 	 1'b0
;    4214		:	dataRd	 = 	 1'b0
;    4215		:	dataRd	 = 	 1'b0
;    4216		:	dataRd	 = 	 1'b0
;    4217		:	dataRd	 = 	 1'b0
;    4218		:	dataRd	 = 	 1'b1
;    4219		:	dataRd	 = 	 1'b0
;    4220		:	dataRd	 = 	 1'b0
;    4221		:	dataRd	 = 	 1'b0
;    4222		:	dataRd	 = 	 1'b0
;    4223		:	dataRd	 = 	 1'b0
;    4224		:	dataRd	 = 	 1'b0
;    4225		:	dataRd	 = 	 1'b0
;    4226		:	dataRd	 = 	 1'b0
;    4227		:	dataRd	 = 	 1'b0
;    4228		:	dataRd	 = 	 1'b0
;    4229		:	dataRd	 = 	 1'b0
;    4230		:	dataRd	 = 	 1'b0
;    4231		:	dataRd	 = 	 1'b0
;    4232		:	dataRd	 = 	 1'b0
;    4233		:	dataRd	 = 	 1'b0
;    4234		:	dataRd	 = 	 1'b1
;    4235		:	dataRd	 = 	 1'b0
;    4236		:	dataRd	 = 	 1'b0
;    4237		:	dataRd	 = 	 1'b0
;    4238		:	dataRd	 = 	 1'b0
;    4239		:	dataRd	 = 	 1'b0
;    4240		:	dataRd	 = 	 1'b0
;    4241		:	dataRd	 = 	 1'b0
;    4242		:	dataRd	 = 	 1'b0
;    4243		:	dataRd	 = 	 1'b0
;    4244		:	dataRd	 = 	 1'b0
;    4245		:	dataRd	 = 	 1'b0
;    4246		:	dataRd	 = 	 1'b0
;    4247		:	dataRd	 = 	 1'b0
;    4248		:	dataRd	 = 	 1'b0
;    4249		:	dataRd	 = 	 1'b0
;    4250		:	dataRd	 = 	 1'b1
;    4251		:	dataRd	 = 	 1'b0
;    4252		:	dataRd	 = 	 1'b0
;    4253		:	dataRd	 = 	 1'b0
;    4254		:	dataRd	 = 	 1'b0
;    4255		:	dataRd	 = 	 1'b0
;    4256		:	dataRd	 = 	 1'b0
;    4257		:	dataRd	 = 	 1'b0
;    4258		:	dataRd	 = 	 1'b0
;    4259		:	dataRd	 = 	 1'b0
;    4260		:	dataRd	 = 	 1'b0
;    4261		:	dataRd	 = 	 1'b0
;    4262		:	dataRd	 = 	 1'b0
;    4263		:	dataRd	 = 	 1'b0
;    4264		:	dataRd	 = 	 1'b0
;    4265		:	dataRd	 = 	 1'b0
;    4266		:	dataRd	 = 	 1'b1
;    4267		:	dataRd	 = 	 1'b0
;    4268		:	dataRd	 = 	 1'b0
;    4269		:	dataRd	 = 	 1'b0
;    4270		:	dataRd	 = 	 1'b0
;    4271		:	dataRd	 = 	 1'b0
;    4272		:	dataRd	 = 	 1'b0
;    4273		:	dataRd	 = 	 1'b0
;    4274		:	dataRd	 = 	 1'b0
;    4275		:	dataRd	 = 	 1'b0
;    4276		:	dataRd	 = 	 1'b0
;    4277		:	dataRd	 = 	 1'b0
;    4278		:	dataRd	 = 	 1'b0
;    4279		:	dataRd	 = 	 1'b0
;    4280		:	dataRd	 = 	 1'b0
;    4281		:	dataRd	 = 	 1'b0
;    4282		:	dataRd	 = 	 1'b1
;    4283		:	dataRd	 = 	 1'b0
;    4284		:	dataRd	 = 	 1'b0
;    4285		:	dataRd	 = 	 1'b0
;    4286		:	dataRd	 = 	 1'b0
;    4287		:	dataRd	 = 	 1'b0
;    4288		:	dataRd	 = 	 1'b0
;    4289		:	dataRd	 = 	 1'b0
;    4290		:	dataRd	 = 	 1'b0
;    4291		:	dataRd	 = 	 1'b0
;    4292		:	dataRd	 = 	 1'b0
;    4293		:	dataRd	 = 	 1'b0
;    4294		:	dataRd	 = 	 1'b0
;    4295		:	dataRd	 = 	 1'b0
;    4296		:	dataRd	 = 	 1'b0
;    4297		:	dataRd	 = 	 1'b0
;    4298		:	dataRd	 = 	 1'b1
;    4299		:	dataRd	 = 	 1'b0
;    4300		:	dataRd	 = 	 1'b0
;    4301		:	dataRd	 = 	 1'b0
;    4302		:	dataRd	 = 	 1'b0
;    4303		:	dataRd	 = 	 1'b0
;    4304		:	dataRd	 = 	 1'b0
;    4305		:	dataRd	 = 	 1'b0
;    4306		:	dataRd	 = 	 1'b0
;    4307		:	dataRd	 = 	 1'b0
;    4308		:	dataRd	 = 	 1'b0
;    4309		:	dataRd	 = 	 1'b0
;    4310		:	dataRd	 = 	 1'b0
;    4311		:	dataRd	 = 	 1'b0
;    4312		:	dataRd	 = 	 1'b0
;    4313		:	dataRd	 = 	 1'b0
;    4314		:	dataRd	 = 	 1'b1
;    4315		:	dataRd	 = 	 1'b0
;    4316		:	dataRd	 = 	 1'b0
;    4317		:	dataRd	 = 	 1'b0
;    4318		:	dataRd	 = 	 1'b0
;    4319		:	dataRd	 = 	 1'b0
;    4320		:	dataRd	 = 	 1'b0
;    4321		:	dataRd	 = 	 1'b0
;    4322		:	dataRd	 = 	 1'b0
;    4323		:	dataRd	 = 	 1'b0
;    4324		:	dataRd	 = 	 1'b0
;    4325		:	dataRd	 = 	 1'b0
;    4326		:	dataRd	 = 	 1'b0
;    4327		:	dataRd	 = 	 1'b0
;    4328		:	dataRd	 = 	 1'b0
;    4329		:	dataRd	 = 	 1'b0
;    4330		:	dataRd	 = 	 1'b1
;    4331		:	dataRd	 = 	 1'b0
;    4332		:	dataRd	 = 	 1'b0
;    4333		:	dataRd	 = 	 1'b0
;    4334		:	dataRd	 = 	 1'b0
;    4335		:	dataRd	 = 	 1'b0
;    4336		:	dataRd	 = 	 1'b0
;    4337		:	dataRd	 = 	 1'b0
;    4338		:	dataRd	 = 	 1'b0
;    4339		:	dataRd	 = 	 1'b0
;    4340		:	dataRd	 = 	 1'b0
;    4341		:	dataRd	 = 	 1'b0
;    4342		:	dataRd	 = 	 1'b0
;    4343		:	dataRd	 = 	 1'b0
;    4344		:	dataRd	 = 	 1'b0
;    4345		:	dataRd	 = 	 1'b0
;    4346		:	dataRd	 = 	 1'b1
;    4347		:	dataRd	 = 	 1'b0
;    4348		:	dataRd	 = 	 1'b0
;    4349		:	dataRd	 = 	 1'b0
;    4350		:	dataRd	 = 	 1'b0
;    4351		:	dataRd	 = 	 1'b0
;    4352		:	dataRd	 = 	 1'b0
;    4353		:	dataRd	 = 	 1'b0
;    4354		:	dataRd	 = 	 1'b0
;    4355		:	dataRd	 = 	 1'b0
;    4356		:	dataRd	 = 	 1'b0
;    4357		:	dataRd	 = 	 1'b0
;    4358		:	dataRd	 = 	 1'b0
;    4359		:	dataRd	 = 	 1'b0
;    4360		:	dataRd	 = 	 1'b0
;    4361		:	dataRd	 = 	 1'b0
;    4362		:	dataRd	 = 	 1'b1
;    4363		:	dataRd	 = 	 1'b0
;    4364		:	dataRd	 = 	 1'b0
;    4365		:	dataRd	 = 	 1'b0
;    4366		:	dataRd	 = 	 1'b0
;    4367		:	dataRd	 = 	 1'b0
;    4368		:	dataRd	 = 	 1'b0
;    4369		:	dataRd	 = 	 1'b0
;    4370		:	dataRd	 = 	 1'b0
;    4371		:	dataRd	 = 	 1'b0
;    4372		:	dataRd	 = 	 1'b0
;    4373		:	dataRd	 = 	 1'b0
;    4374		:	dataRd	 = 	 1'b0
;    4375		:	dataRd	 = 	 1'b0
;    4376		:	dataRd	 = 	 1'b0
;    4377		:	dataRd	 = 	 1'b0
;    4378		:	dataRd	 = 	 1'b1
;    4379		:	dataRd	 = 	 1'b0
;    4380		:	dataRd	 = 	 1'b0
;    4381		:	dataRd	 = 	 1'b0
;    4382		:	dataRd	 = 	 1'b0
;    4383		:	dataRd	 = 	 1'b0
;    4384		:	dataRd	 = 	 1'b0
;    4385		:	dataRd	 = 	 1'b0
;    4386		:	dataRd	 = 	 1'b0
;    4387		:	dataRd	 = 	 1'b0
;    4388		:	dataRd	 = 	 1'b0
;    4389		:	dataRd	 = 	 1'b0
;    4390		:	dataRd	 = 	 1'b0
;    4391		:	dataRd	 = 	 1'b0
;    4392		:	dataRd	 = 	 1'b0
;    4393		:	dataRd	 = 	 1'b0
;    4394		:	dataRd	 = 	 1'b1
;    4395		:	dataRd	 = 	 1'b0
;    4396		:	dataRd	 = 	 1'b0
;    4397		:	dataRd	 = 	 1'b0
;    4398		:	dataRd	 = 	 1'b0
;    4399		:	dataRd	 = 	 1'b0
;    4400		:	dataRd	 = 	 1'b0
;    4401		:	dataRd	 = 	 1'b0
;    4402		:	dataRd	 = 	 1'b0
;    4403		:	dataRd	 = 	 1'b0
;    4404		:	dataRd	 = 	 1'b0
;    4405		:	dataRd	 = 	 1'b0
;    4406		:	dataRd	 = 	 1'b0
;    4407		:	dataRd	 = 	 1'b0
;    4408		:	dataRd	 = 	 1'b0
;    4409		:	dataRd	 = 	 1'b0
;    4410		:	dataRd	 = 	 1'b1
;    4411		:	dataRd	 = 	 1'b0
;    4412		:	dataRd	 = 	 1'b0
;    4413		:	dataRd	 = 	 1'b0
;    4414		:	dataRd	 = 	 1'b0
;    4415		:	dataRd	 = 	 1'b0
;    4416		:	dataRd	 = 	 1'b0
;    4417		:	dataRd	 = 	 1'b0
;    4418		:	dataRd	 = 	 1'b0
;    4419		:	dataRd	 = 	 1'b0
;    4420		:	dataRd	 = 	 1'b0
;    4421		:	dataRd	 = 	 1'b0
;    4422		:	dataRd	 = 	 1'b0
;    4423		:	dataRd	 = 	 1'b0
;    4424		:	dataRd	 = 	 1'b0
;    4425		:	dataRd	 = 	 1'b0
;    4426		:	dataRd	 = 	 1'b1
;    4427		:	dataRd	 = 	 1'b0
;    4428		:	dataRd	 = 	 1'b0
;    4429		:	dataRd	 = 	 1'b0
;    4430		:	dataRd	 = 	 1'b0
;    4431		:	dataRd	 = 	 1'b0
;    4432		:	dataRd	 = 	 1'b0
;    4433		:	dataRd	 = 	 1'b0
;    4434		:	dataRd	 = 	 1'b0
;    4435		:	dataRd	 = 	 1'b0
;    4436		:	dataRd	 = 	 1'b0
;    4437		:	dataRd	 = 	 1'b0
;    4438		:	dataRd	 = 	 1'b0
;    4439		:	dataRd	 = 	 1'b0
;    4440		:	dataRd	 = 	 1'b0
;    4441		:	dataRd	 = 	 1'b0
;    4442		:	dataRd	 = 	 1'b0
;    4443		:	dataRd	 = 	 1'b1
;    4444		:	dataRd	 = 	 1'b0
;    4445		:	dataRd	 = 	 1'b0
;    4446		:	dataRd	 = 	 1'b0
;    4447		:	dataRd	 = 	 1'b0
;    4448		:	dataRd	 = 	 1'b0
;    4449		:	dataRd	 = 	 1'b0
;    4450		:	dataRd	 = 	 1'b0
;    4451		:	dataRd	 = 	 1'b0
;    4452		:	dataRd	 = 	 1'b0
;    4453		:	dataRd	 = 	 1'b0
;    4454		:	dataRd	 = 	 1'b0
;    4455		:	dataRd	 = 	 1'b0
;    4456		:	dataRd	 = 	 1'b0
;    4457		:	dataRd	 = 	 1'b0
;    4458		:	dataRd	 = 	 1'b0
;    4459		:	dataRd	 = 	 1'b0
;    4460		:	dataRd	 = 	 1'b0
;    4461		:	dataRd	 = 	 1'b0
;    4462		:	dataRd	 = 	 1'b0
;    4463		:	dataRd	 = 	 1'b0
;    4464		:	dataRd	 = 	 1'b0
;    4465		:	dataRd	 = 	 1'b0
;    4466		:	dataRd	 = 	 1'b0
;    4467		:	dataRd	 = 	 1'b0
;    4468		:	dataRd	 = 	 1'b0
;    4469		:	dataRd	 = 	 1'b0
;    4470		:	dataRd	 = 	 1'b0
;    4471		:	dataRd	 = 	 1'b0
;    4472		:	dataRd	 = 	 1'b0
;    4473		:	dataRd	 = 	 1'b0
;    4474		:	dataRd	 = 	 1'b0
;    4475		:	dataRd	 = 	 1'b0
;    4476		:	dataRd	 = 	 1'b0
;    4477		:	dataRd	 = 	 1'b0
;    4478		:	dataRd	 = 	 1'b0
;    4479		:	dataRd	 = 	 1'b0
;    4480		:	dataRd	 = 	 1'b0
;    4481		:	dataRd	 = 	 1'b0
;    4482		:	dataRd	 = 	 1'b0
;    4483		:	dataRd	 = 	 1'b0
;    4484		:	dataRd	 = 	 1'b0
;    4485		:	dataRd	 = 	 1'b1
;    4486		:	dataRd	 = 	 1'b1
;    4487		:	dataRd	 = 	 1'b1
;    4488		:	dataRd	 = 	 1'b1
;    4489		:	dataRd	 = 	 1'b1
;    4490		:	dataRd	 = 	 1'b1
;    4491		:	dataRd	 = 	 1'b1
;    4492		:	dataRd	 = 	 1'b1
;    4493		:	dataRd	 = 	 1'b0
;    4494		:	dataRd	 = 	 1'b0
;    4495		:	dataRd	 = 	 1'b0
;    4496		:	dataRd	 = 	 1'b0
;    4497		:	dataRd	 = 	 1'b0
;    4498		:	dataRd	 = 	 1'b0
;    4499		:	dataRd	 = 	 1'b0
;    4500		:	dataRd	 = 	 1'b0
;    4501		:	dataRd	 = 	 1'b1
;    4502		:	dataRd	 = 	 1'b1
;    4503		:	dataRd	 = 	 1'b1
;    4504		:	dataRd	 = 	 1'b1
;    4505		:	dataRd	 = 	 1'b1
;    4506		:	dataRd	 = 	 1'b1
;    4507		:	dataRd	 = 	 1'b1
;    4508		:	dataRd	 = 	 1'b1
;    4509		:	dataRd	 = 	 1'b1
;    4510		:	dataRd	 = 	 1'b0
;    4511		:	dataRd	 = 	 1'b0
;    4512		:	dataRd	 = 	 1'b0
;    4513		:	dataRd	 = 	 1'b0
;    4514		:	dataRd	 = 	 1'b0
;    4515		:	dataRd	 = 	 1'b0
;    4516		:	dataRd	 = 	 1'b0
;    4517		:	dataRd	 = 	 1'b0
;    4518		:	dataRd	 = 	 1'b0
;    4519		:	dataRd	 = 	 1'b0
;    4520		:	dataRd	 = 	 1'b0
;    4521		:	dataRd	 = 	 1'b0
;    4522		:	dataRd	 = 	 1'b0
;    4523		:	dataRd	 = 	 1'b0
;    4524		:	dataRd	 = 	 1'b0
;    4525		:	dataRd	 = 	 1'b0
;    4526		:	dataRd	 = 	 1'b0
;    4527		:	dataRd	 = 	 1'b0
;    4528		:	dataRd	 = 	 1'b0
;    4529		:	dataRd	 = 	 1'b0
;    4530		:	dataRd	 = 	 1'b0
;    4531		:	dataRd	 = 	 1'b0
;    4532		:	dataRd	 = 	 1'b0
;    4533		:	dataRd	 = 	 1'b0
;    4534		:	dataRd	 = 	 1'b0
;    4535		:	dataRd	 = 	 1'b0
;    4536		:	dataRd	 = 	 1'b0
;    4537		:	dataRd	 = 	 1'b0
;    4538		:	dataRd	 = 	 1'b0
;    4539		:	dataRd	 = 	 1'b0
;    4540		:	dataRd	 = 	 1'b0
;    4541		:	dataRd	 = 	 1'b0
;    4542		:	dataRd	 = 	 1'b0
;    4543		:	dataRd	 = 	 1'b0
;    4544		:	dataRd	 = 	 1'b0
;    4545		:	dataRd	 = 	 1'b0
;    4546		:	dataRd	 = 	 1'b0
;    4547		:	dataRd	 = 	 1'b0
;    4548		:	dataRd	 = 	 1'b0
;    4549		:	dataRd	 = 	 1'b0
;    4550		:	dataRd	 = 	 1'b0
;    4551		:	dataRd	 = 	 1'b0
;    4552		:	dataRd	 = 	 1'b0
;    4553		:	dataRd	 = 	 1'b0
;    4554		:	dataRd	 = 	 1'b0
;    4555		:	dataRd	 = 	 1'b0
;    4556		:	dataRd	 = 	 1'b0
;    4557		:	dataRd	 = 	 1'b0
;    4558		:	dataRd	 = 	 1'b0
;    4559		:	dataRd	 = 	 1'b0
;    4560		:	dataRd	 = 	 1'b0
;    4561		:	dataRd	 = 	 1'b0
;    4562		:	dataRd	 = 	 1'b0
;    4563		:	dataRd	 = 	 1'b0
;    4564		:	dataRd	 = 	 1'b0
;    4565		:	dataRd	 = 	 1'b0
;    4566		:	dataRd	 = 	 1'b0
;    4567		:	dataRd	 = 	 1'b0
;    4568		:	dataRd	 = 	 1'b0
;    4569		:	dataRd	 = 	 1'b0
;    4570		:	dataRd	 = 	 1'b0
;    4571		:	dataRd	 = 	 1'b0
;    4572		:	dataRd	 = 	 1'b0
;    4573		:	dataRd	 = 	 1'b0
;    4574		:	dataRd	 = 	 1'b0
;    4575		:	dataRd	 = 	 1'b0
;    4576		:	dataRd	 = 	 1'b1
;    4577		:	dataRd	 = 	 1'b0
;    4578		:	dataRd	 = 	 1'b0
;    4579		:	dataRd	 = 	 1'b0
;    4580		:	dataRd	 = 	 1'b0
;    4581		:	dataRd	 = 	 1'b0
;    4582		:	dataRd	 = 	 1'b0
;    4583		:	dataRd	 = 	 1'b0
;    4584		:	dataRd	 = 	 1'b0
;    4585		:	dataRd	 = 	 1'b0
;    4586		:	dataRd	 = 	 1'b0
;    4587		:	dataRd	 = 	 1'b0
;    4588		:	dataRd	 = 	 1'b0
;    4589		:	dataRd	 = 	 1'b0
;    4590		:	dataRd	 = 	 1'b0
;    4591		:	dataRd	 = 	 1'b0
;    4592		:	dataRd	 = 	 1'b0
;    4593		:	dataRd	 = 	 1'b0
;    4594		:	dataRd	 = 	 1'b0
;    4595		:	dataRd	 = 	 1'b0
;    4596		:	dataRd	 = 	 1'b0
;    4597		:	dataRd	 = 	 1'b0
;    4598		:	dataRd	 = 	 1'b0
;    4599		:	dataRd	 = 	 1'b0
;    4600		:	dataRd	 = 	 1'b0
;    4601		:	dataRd	 = 	 1'b0
;    4602		:	dataRd	 = 	 1'b0
;    4603		:	dataRd	 = 	 1'b0
;    4604		:	dataRd	 = 	 1'b0
;    4605		:	dataRd	 = 	 1'b0
;    4606		:	dataRd	 = 	 1'b0
;    4607		:	dataRd	 = 	 1'b0
;    4608		:	dataRd	 = 	 1'b0
;    4609		:	dataRd	 = 	 1'b0
;    4610		:	dataRd	 = 	 1'b0
;    4611		:	dataRd	 = 	 1'b0
;    4612		:	dataRd	 = 	 1'b0
;    4613		:	dataRd	 = 	 1'b0
;    4614		:	dataRd	 = 	 1'b0
;    4615		:	dataRd	 = 	 1'b0
;    4616		:	dataRd	 = 	 1'b0
;    4617		:	dataRd	 = 	 1'b0
;    4618		:	dataRd	 = 	 1'b0
;    4619		:	dataRd	 = 	 1'b0
;    4620		:	dataRd	 = 	 1'b0
;    4621		:	dataRd	 = 	 1'b0
;    4622		:	dataRd	 = 	 1'b0
;    4623		:	dataRd	 = 	 1'b0
;    4624		:	dataRd	 = 	 1'b0
;    4625		:	dataRd	 = 	 1'b0
;    4626		:	dataRd	 = 	 1'b0
;    4627		:	dataRd	 = 	 1'b0
;    4628		:	dataRd	 = 	 1'b0
;    4629		:	dataRd	 = 	 1'b0
;    4630		:	dataRd	 = 	 1'b0
;    4631		:	dataRd	 = 	 1'b0
;    4632		:	dataRd	 = 	 1'b0
;    4633		:	dataRd	 = 	 1'b0
;    4634		:	dataRd	 = 	 1'b0
;    4635		:	dataRd	 = 	 1'b0
;    4636		:	dataRd	 = 	 1'b0
;    4637		:	dataRd	 = 	 1'b0
;    4638		:	dataRd	 = 	 1'b0
;    4639		:	dataRd	 = 	 1'b0
;    4640		:	dataRd	 = 	 1'b0
;    4641		:	dataRd	 = 	 1'b0
;    4642		:	dataRd	 = 	 1'b0
;    4643		:	dataRd	 = 	 1'b1
;    4644		:	dataRd	 = 	 1'b0
;    4645		:	dataRd	 = 	 1'b0
;    4646		:	dataRd	 = 	 1'b0
;    4647		:	dataRd	 = 	 1'b0
;    4648		:	dataRd	 = 	 1'b0
;    4649		:	dataRd	 = 	 1'b0
;    4650		:	dataRd	 = 	 1'b0
;    4651		:	dataRd	 = 	 1'b0
;    4652		:	dataRd	 = 	 1'b0
;    4653		:	dataRd	 = 	 1'b0
;    4654		:	dataRd	 = 	 1'b0
;    4655		:	dataRd	 = 	 1'b0
;    4656		:	dataRd	 = 	 1'b0
;    4657		:	dataRd	 = 	 1'b0
;    4658		:	dataRd	 = 	 1'b0
;    4659		:	dataRd	 = 	 1'b0
;    4660		:	dataRd	 = 	 1'b0
;    4661		:	dataRd	 = 	 1'b0
;    4662		:	dataRd	 = 	 1'b0
;    4663		:	dataRd	 = 	 1'b0
;    4664		:	dataRd	 = 	 1'b0
;    4665		:	dataRd	 = 	 1'b0
;    4666		:	dataRd	 = 	 1'b0
;    4667		:	dataRd	 = 	 1'b0
;    4668		:	dataRd	 = 	 1'b0
;    4669		:	dataRd	 = 	 1'b0
;    4670		:	dataRd	 = 	 1'b0
;    4671		:	dataRd	 = 	 1'b0
;    4672		:	dataRd	 = 	 1'b0
;    4673		:	dataRd	 = 	 1'b0
;    4674		:	dataRd	 = 	 1'b0
;    4675		:	dataRd	 = 	 1'b0
;    4676		:	dataRd	 = 	 1'b0
;    4677		:	dataRd	 = 	 1'b0
;    4678		:	dataRd	 = 	 1'b0
;    4679		:	dataRd	 = 	 1'b0
;    4680		:	dataRd	 = 	 1'b0
;    4681		:	dataRd	 = 	 1'b0
;    4682		:	dataRd	 = 	 1'b0
;    4683		:	dataRd	 = 	 1'b0
;    4684		:	dataRd	 = 	 1'b0
;    4685		:	dataRd	 = 	 1'b0
;    4686		:	dataRd	 = 	 1'b0
;    4687		:	dataRd	 = 	 1'b0
;    4688		:	dataRd	 = 	 1'b0
;    4689		:	dataRd	 = 	 1'b0
;    4690		:	dataRd	 = 	 1'b0
;    4691		:	dataRd	 = 	 1'b0
;    4692		:	dataRd	 = 	 1'b0
;    4693		:	dataRd	 = 	 1'b0
;    4694		:	dataRd	 = 	 1'b0
;    4695		:	dataRd	 = 	 1'b0
;    4696		:	dataRd	 = 	 1'b0
;    4697		:	dataRd	 = 	 1'b0
;    4698		:	dataRd	 = 	 1'b0
;    4699		:	dataRd	 = 	 1'b0
;    4700		:	dataRd	 = 	 1'b0
;    4701		:	dataRd	 = 	 1'b0
;    4702		:	dataRd	 = 	 1'b0
;    4703		:	dataRd	 = 	 1'b0
;    4704		:	dataRd	 = 	 1'b0
;    4705		:	dataRd	 = 	 1'b0
;    4706		:	dataRd	 = 	 1'b0
;    4707		:	dataRd	 = 	 1'b0
;    4708		:	dataRd	 = 	 1'b0
;    4709		:	dataRd	 = 	 1'b0
;    4710		:	dataRd	 = 	 1'b1
;    4711		:	dataRd	 = 	 1'b0
;    4712		:	dataRd	 = 	 1'b0
;    4713		:	dataRd	 = 	 1'b0
;    4714		:	dataRd	 = 	 1'b0
;    4715		:	dataRd	 = 	 1'b0
;    4716		:	dataRd	 = 	 1'b0
;    4717		:	dataRd	 = 	 1'b0
;    4718		:	dataRd	 = 	 1'b0
;    4719		:	dataRd	 = 	 1'b0
;    4720		:	dataRd	 = 	 1'b0
;    4721		:	dataRd	 = 	 1'b0
;    4722		:	dataRd	 = 	 1'b0
;    4723		:	dataRd	 = 	 1'b0
;    4724		:	dataRd	 = 	 1'b0
;    4725		:	dataRd	 = 	 1'b0
;    4726		:	dataRd	 = 	 1'b0
;    4727		:	dataRd	 = 	 1'b0
;    4728		:	dataRd	 = 	 1'b0
;    4729		:	dataRd	 = 	 1'b0
;    4730		:	dataRd	 = 	 1'b0
;    4731		:	dataRd	 = 	 1'b0
;    4732		:	dataRd	 = 	 1'b0
;    4733		:	dataRd	 = 	 1'b0
;    4734		:	dataRd	 = 	 1'b0
;    4735		:	dataRd	 = 	 1'b0
;    4736		:	dataRd	 = 	 1'b0
;    4737		:	dataRd	 = 	 1'b0
;    4738		:	dataRd	 = 	 1'b0
;    4739		:	dataRd	 = 	 1'b0
;    4740		:	dataRd	 = 	 1'b0
;    4741		:	dataRd	 = 	 1'b0
;    4742		:	dataRd	 = 	 1'b0
;    4743		:	dataRd	 = 	 1'b0
;    4744		:	dataRd	 = 	 1'b0
;    4745		:	dataRd	 = 	 1'b0
;    4746		:	dataRd	 = 	 1'b0
;    4747		:	dataRd	 = 	 1'b0
;    4748		:	dataRd	 = 	 1'b0
;    4749		:	dataRd	 = 	 1'b0
;    4750		:	dataRd	 = 	 1'b0
;    4751		:	dataRd	 = 	 1'b0
;    4752		:	dataRd	 = 	 1'b0
;    4753		:	dataRd	 = 	 1'b0
;    4754		:	dataRd	 = 	 1'b0
;    4755		:	dataRd	 = 	 1'b0
;    4756		:	dataRd	 = 	 1'b0
;    4757		:	dataRd	 = 	 1'b0
;    4758		:	dataRd	 = 	 1'b0
;    4759		:	dataRd	 = 	 1'b0
;    4760		:	dataRd	 = 	 1'b0
;    4761		:	dataRd	 = 	 1'b0
;    4762		:	dataRd	 = 	 1'b0
;    4763		:	dataRd	 = 	 1'b0
;    4764		:	dataRd	 = 	 1'b0
;    4765		:	dataRd	 = 	 1'b0
;    4766		:	dataRd	 = 	 1'b0
;    4767		:	dataRd	 = 	 1'b0
;    4768		:	dataRd	 = 	 1'b0
;    4769		:	dataRd	 = 	 1'b0
;    4770		:	dataRd	 = 	 1'b0
;    4771		:	dataRd	 = 	 1'b0
;    4772		:	dataRd	 = 	 1'b0
;    4773		:	dataRd	 = 	 1'b0
;    4774		:	dataRd	 = 	 1'b0
;    4775		:	dataRd	 = 	 1'b0
;    4776		:	dataRd	 = 	 1'b0
;    4777		:	dataRd	 = 	 1'b1
;    4778		:	dataRd	 = 	 1'b0
;    4779		:	dataRd	 = 	 1'b0
;    4780		:	dataRd	 = 	 1'b0
;    4781		:	dataRd	 = 	 1'b0
;    4782		:	dataRd	 = 	 1'b0
;    4783		:	dataRd	 = 	 1'b0
;    4784		:	dataRd	 = 	 1'b0
;    4785		:	dataRd	 = 	 1'b0
;    4786		:	dataRd	 = 	 1'b0
;    4787		:	dataRd	 = 	 1'b0
;    4788		:	dataRd	 = 	 1'b0
;    4789		:	dataRd	 = 	 1'b0
;    4790		:	dataRd	 = 	 1'b0
;    4791		:	dataRd	 = 	 1'b0
;    4792		:	dataRd	 = 	 1'b0
;    4793		:	dataRd	 = 	 1'b0
;    4794		:	dataRd	 = 	 1'b0
;    4795		:	dataRd	 = 	 1'b0
;    4796		:	dataRd	 = 	 1'b0
;    4797		:	dataRd	 = 	 1'b0
;    4798		:	dataRd	 = 	 1'b0
;    4799		:	dataRd	 = 	 1'b0
;    4800		:	dataRd	 = 	 1'b0
;    4801		:	dataRd	 = 	 1'b0
;    4802		:	dataRd	 = 	 1'b0
;    4803		:	dataRd	 = 	 1'b0
;    4804		:	dataRd	 = 	 1'b0
;    4805		:	dataRd	 = 	 1'b0
;    4806		:	dataRd	 = 	 1'b0
;    4807		:	dataRd	 = 	 1'b0
;    4808		:	dataRd	 = 	 1'b0
;    4809		:	dataRd	 = 	 1'b0
;    4810		:	dataRd	 = 	 1'b0
;    4811		:	dataRd	 = 	 1'b0
;    4812		:	dataRd	 = 	 1'b0
;    4813		:	dataRd	 = 	 1'b0
;    4814		:	dataRd	 = 	 1'b0
;    4815		:	dataRd	 = 	 1'b0
;    4816		:	dataRd	 = 	 1'b0
;    4817		:	dataRd	 = 	 1'b0
;    4818		:	dataRd	 = 	 1'b0
;    4819		:	dataRd	 = 	 1'b0
;    4820		:	dataRd	 = 	 1'b0
;    4821		:	dataRd	 = 	 1'b0
;    4822		:	dataRd	 = 	 1'b0
;    4823		:	dataRd	 = 	 1'b0
;    4824		:	dataRd	 = 	 1'b0
;    4825		:	dataRd	 = 	 1'b0
;    4826		:	dataRd	 = 	 1'b0
;    4827		:	dataRd	 = 	 1'b0
;    4828		:	dataRd	 = 	 1'b0
;    4829		:	dataRd	 = 	 1'b0
;    4830		:	dataRd	 = 	 1'b0
;    4831		:	dataRd	 = 	 1'b0
;    4832		:	dataRd	 = 	 1'b0
;    4833		:	dataRd	 = 	 1'b0
;    4834		:	dataRd	 = 	 1'b0
;    4835		:	dataRd	 = 	 1'b0
;    4836		:	dataRd	 = 	 1'b0
;    4837		:	dataRd	 = 	 1'b0
;    4838		:	dataRd	 = 	 1'b0
;    4839		:	dataRd	 = 	 1'b0
;    4840		:	dataRd	 = 	 1'b0
;    4841		:	dataRd	 = 	 1'b0
;    4842		:	dataRd	 = 	 1'b0
;    4843		:	dataRd	 = 	 1'b0
;    4844		:	dataRd	 = 	 1'b1
;    4845		:	dataRd	 = 	 1'b0
;    4846		:	dataRd	 = 	 1'b0
;    4847		:	dataRd	 = 	 1'b0
;    4848		:	dataRd	 = 	 1'b0
;    4849		:	dataRd	 = 	 1'b0
;    4850		:	dataRd	 = 	 1'b0
;    4851		:	dataRd	 = 	 1'b0
;    4852		:	dataRd	 = 	 1'b0
;    4853		:	dataRd	 = 	 1'b0
;    4854		:	dataRd	 = 	 1'b0
;    4855		:	dataRd	 = 	 1'b0
;    4856		:	dataRd	 = 	 1'b0
;    4857		:	dataRd	 = 	 1'b0
;    4858		:	dataRd	 = 	 1'b0
;    4859		:	dataRd	 = 	 1'b0
;    4860		:	dataRd	 = 	 1'b0
;    4861		:	dataRd	 = 	 1'b0
;    4862		:	dataRd	 = 	 1'b0
;    4863		:	dataRd	 = 	 1'b0
;    4864		:	dataRd	 = 	 1'b0
;    4865		:	dataRd	 = 	 1'b0
;    4866		:	dataRd	 = 	 1'b0
;    4867		:	dataRd	 = 	 1'b0
;    4868		:	dataRd	 = 	 1'b0
;    4869		:	dataRd	 = 	 1'b0
;    4870		:	dataRd	 = 	 1'b0
;    4871		:	dataRd	 = 	 1'b0
;    4872		:	dataRd	 = 	 1'b0
;    4873		:	dataRd	 = 	 1'b0
;    4874		:	dataRd	 = 	 1'b0
;    4875		:	dataRd	 = 	 1'b0
;    4876		:	dataRd	 = 	 1'b0
;    4877		:	dataRd	 = 	 1'b0
;    4878		:	dataRd	 = 	 1'b0
;    4879		:	dataRd	 = 	 1'b0
;    4880		:	dataRd	 = 	 1'b0
;    4881		:	dataRd	 = 	 1'b0
;    4882		:	dataRd	 = 	 1'b0
;    4883		:	dataRd	 = 	 1'b0
;    4884		:	dataRd	 = 	 1'b0
;    4885		:	dataRd	 = 	 1'b0
;    4886		:	dataRd	 = 	 1'b0
;    4887		:	dataRd	 = 	 1'b0
;    4888		:	dataRd	 = 	 1'b0
;    4889		:	dataRd	 = 	 1'b0
;    4890		:	dataRd	 = 	 1'b0
;    4891		:	dataRd	 = 	 1'b0
;    4892		:	dataRd	 = 	 1'b0
;    4893		:	dataRd	 = 	 1'b0
;    4894		:	dataRd	 = 	 1'b0
;    4895		:	dataRd	 = 	 1'b0
;    4896		:	dataRd	 = 	 1'b0
;    4897		:	dataRd	 = 	 1'b0
;    4898		:	dataRd	 = 	 1'b0
;    4899		:	dataRd	 = 	 1'b0
;    4900		:	dataRd	 = 	 1'b0
;    4901		:	dataRd	 = 	 1'b0
;    4902		:	dataRd	 = 	 1'b0
;    4903		:	dataRd	 = 	 1'b0
;    4904		:	dataRd	 = 	 1'b0
;    4905		:	dataRd	 = 	 1'b0
;    4906		:	dataRd	 = 	 1'b0
;    4907		:	dataRd	 = 	 1'b0
;    4908		:	dataRd	 = 	 1'b0
;    4909		:	dataRd	 = 	 1'b0
;    4910		:	dataRd	 = 	 1'b0
;    4911		:	dataRd	 = 	 1'b1
;    4912		:	dataRd	 = 	 1'b0
;    4913		:	dataRd	 = 	 1'b0
;    4914		:	dataRd	 = 	 1'b0
;    4915		:	dataRd	 = 	 1'b0
;    4916		:	dataRd	 = 	 1'b0
;    4917		:	dataRd	 = 	 1'b0
;    4918		:	dataRd	 = 	 1'b0
;    4919		:	dataRd	 = 	 1'b0
;    4920		:	dataRd	 = 	 1'b0
;    4921		:	dataRd	 = 	 1'b0
;    4922		:	dataRd	 = 	 1'b0
;    4923		:	dataRd	 = 	 1'b0
;    4924		:	dataRd	 = 	 1'b0
;    4925		:	dataRd	 = 	 1'b0
;    4926		:	dataRd	 = 	 1'b0
;    4927		:	dataRd	 = 	 1'b0
;    4928		:	dataRd	 = 	 1'b0
;    4929		:	dataRd	 = 	 1'b0
;    4930		:	dataRd	 = 	 1'b0
;    4931		:	dataRd	 = 	 1'b0
;    4932		:	dataRd	 = 	 1'b0
;    4933		:	dataRd	 = 	 1'b0
;    4934		:	dataRd	 = 	 1'b0
;    4935		:	dataRd	 = 	 1'b0
;    4936		:	dataRd	 = 	 1'b0
;    4937		:	dataRd	 = 	 1'b0
;    4938		:	dataRd	 = 	 1'b0
;    4939		:	dataRd	 = 	 1'b0
;    4940		:	dataRd	 = 	 1'b0
;    4941		:	dataRd	 = 	 1'b0
;    4942		:	dataRd	 = 	 1'b0
;    4943		:	dataRd	 = 	 1'b0
;    4944		:	dataRd	 = 	 1'b0
;    4945		:	dataRd	 = 	 1'b0
;    4946		:	dataRd	 = 	 1'b0
;    4947		:	dataRd	 = 	 1'b0
;    4948		:	dataRd	 = 	 1'b0
;    4949		:	dataRd	 = 	 1'b0
;    4950		:	dataRd	 = 	 1'b0
;    4951		:	dataRd	 = 	 1'b0
;    4952		:	dataRd	 = 	 1'b0
;    4953		:	dataRd	 = 	 1'b0
;    4954		:	dataRd	 = 	 1'b0
;    4955		:	dataRd	 = 	 1'b0
;    4956		:	dataRd	 = 	 1'b0
;    4957		:	dataRd	 = 	 1'b0
;    4958		:	dataRd	 = 	 1'b0
;    4959		:	dataRd	 = 	 1'b0
;    4960		:	dataRd	 = 	 1'b0
;    4961		:	dataRd	 = 	 1'b0
;    4962		:	dataRd	 = 	 1'b0
;    4963		:	dataRd	 = 	 1'b0
;    4964		:	dataRd	 = 	 1'b0
;    4965		:	dataRd	 = 	 1'b0
;    4966		:	dataRd	 = 	 1'b0
;    4967		:	dataRd	 = 	 1'b0
;    4968		:	dataRd	 = 	 1'b0
;    4969		:	dataRd	 = 	 1'b0
;    4970		:	dataRd	 = 	 1'b0
;    4971		:	dataRd	 = 	 1'b0
;    4972		:	dataRd	 = 	 1'b0
;    4973		:	dataRd	 = 	 1'b0
;    4974		:	dataRd	 = 	 1'b0
;    4975		:	dataRd	 = 	 1'b0
;    4976		:	dataRd	 = 	 1'b0
;    4977		:	dataRd	 = 	 1'b0
;    4978		:	dataRd	 = 	 1'b1
;    4979		:	dataRd	 = 	 1'b0
;    4980		:	dataRd	 = 	 1'b0
;    4981		:	dataRd	 = 	 1'b0
;    4982		:	dataRd	 = 	 1'b0
;    4983		:	dataRd	 = 	 1'b0
;    4984		:	dataRd	 = 	 1'b0
;    4985		:	dataRd	 = 	 1'b0
;    4986		:	dataRd	 = 	 1'b0
;    4987		:	dataRd	 = 	 1'b0
;    4988		:	dataRd	 = 	 1'b0
;    4989		:	dataRd	 = 	 1'b0
;    4990		:	dataRd	 = 	 1'b0
;    4991		:	dataRd	 = 	 1'b0
;    4992		:	dataRd	 = 	 1'b0
;    4993		:	dataRd	 = 	 1'b0
;    4994		:	dataRd	 = 	 1'b0
;    4995		:	dataRd	 = 	 1'b0
;    4996		:	dataRd	 = 	 1'b0
;    4997		:	dataRd	 = 	 1'b0
;    4998		:	dataRd	 = 	 1'b0
;    4999		:	dataRd	 = 	 1'b0
;    5000		:	dataRd	 = 	 1'b0
;    5001		:	dataRd	 = 	 1'b0
;    5002		:	dataRd	 = 	 1'b0
;    5003		:	dataRd	 = 	 1'b0
;    5004		:	dataRd	 = 	 1'b0
;    5005		:	dataRd	 = 	 1'b0
;    5006		:	dataRd	 = 	 1'b0
;    5007		:	dataRd	 = 	 1'b0
;    5008		:	dataRd	 = 	 1'b0
;    5009		:	dataRd	 = 	 1'b0
;    5010		:	dataRd	 = 	 1'b0
;    5011		:	dataRd	 = 	 1'b0
;    5012		:	dataRd	 = 	 1'b0
;    5013		:	dataRd	 = 	 1'b0
;    5014		:	dataRd	 = 	 1'b0
;    5015		:	dataRd	 = 	 1'b0
;    5016		:	dataRd	 = 	 1'b0
;    5017		:	dataRd	 = 	 1'b0
;    5018		:	dataRd	 = 	 1'b0
;    5019		:	dataRd	 = 	 1'b0
;    5020		:	dataRd	 = 	 1'b0
;    5021		:	dataRd	 = 	 1'b0
;    5022		:	dataRd	 = 	 1'b0
;    5023		:	dataRd	 = 	 1'b0
;    5024		:	dataRd	 = 	 1'b0
;    5025		:	dataRd	 = 	 1'b0
;    5026		:	dataRd	 = 	 1'b0
;    5027		:	dataRd	 = 	 1'b0
;    5028		:	dataRd	 = 	 1'b0
;    5029		:	dataRd	 = 	 1'b0
;    5030		:	dataRd	 = 	 1'b0
;    5031		:	dataRd	 = 	 1'b0
;    5032		:	dataRd	 = 	 1'b0
;    5033		:	dataRd	 = 	 1'b0
;    5034		:	dataRd	 = 	 1'b0
;    5035		:	dataRd	 = 	 1'b0
;    5036		:	dataRd	 = 	 1'b0
;    5037		:	dataRd	 = 	 1'b0
;    5038		:	dataRd	 = 	 1'b0
;    5039		:	dataRd	 = 	 1'b0
;    5040		:	dataRd	 = 	 1'b0
;    5041		:	dataRd	 = 	 1'b0
;    5042		:	dataRd	 = 	 1'b0
;    5043		:	dataRd	 = 	 1'b0
;    5044		:	dataRd	 = 	 1'b0
;    5045		:	dataRd	 = 	 1'b1
;    5046		:	dataRd	 = 	 1'b0
;    5047		:	dataRd	 = 	 1'b0
;    5048		:	dataRd	 = 	 1'b0
;    5049		:	dataRd	 = 	 1'b0
;    5050		:	dataRd	 = 	 1'b0
;    5051		:	dataRd	 = 	 1'b0
;    5052		:	dataRd	 = 	 1'b0
;    5053		:	dataRd	 = 	 1'b0
;    5054		:	dataRd	 = 	 1'b0
;    5055		:	dataRd	 = 	 1'b0
;    5056		:	dataRd	 = 	 1'b0
;    5057		:	dataRd	 = 	 1'b0
;    5058		:	dataRd	 = 	 1'b0
;    5059		:	dataRd	 = 	 1'b0
;    5060		:	dataRd	 = 	 1'b0
;    5061		:	dataRd	 = 	 1'b0
;    5062		:	dataRd	 = 	 1'b0
;    5063		:	dataRd	 = 	 1'b0
;    5064		:	dataRd	 = 	 1'b0
;    5065		:	dataRd	 = 	 1'b0
;    5066		:	dataRd	 = 	 1'b0
;    5067		:	dataRd	 = 	 1'b0
;    5068		:	dataRd	 = 	 1'b0
;    5069		:	dataRd	 = 	 1'b0
;    5070		:	dataRd	 = 	 1'b0
;    5071		:	dataRd	 = 	 1'b0
;    5072		:	dataRd	 = 	 1'b0
;    5073		:	dataRd	 = 	 1'b0
;    5074		:	dataRd	 = 	 1'b0
;    5075		:	dataRd	 = 	 1'b0
;    5076		:	dataRd	 = 	 1'b0
;    5077		:	dataRd	 = 	 1'b0
;    5078		:	dataRd	 = 	 1'b0
;    5079		:	dataRd	 = 	 1'b0
;    5080		:	dataRd	 = 	 1'b0
;    5081		:	dataRd	 = 	 1'b0
;    5082		:	dataRd	 = 	 1'b0
;    5083		:	dataRd	 = 	 1'b0
;    5084		:	dataRd	 = 	 1'b0
;    5085		:	dataRd	 = 	 1'b0
;    5086		:	dataRd	 = 	 1'b0
;    5087		:	dataRd	 = 	 1'b0
;    5088		:	dataRd	 = 	 1'b0
;    5089		:	dataRd	 = 	 1'b0
;    5090		:	dataRd	 = 	 1'b0
;    5091		:	dataRd	 = 	 1'b0
;    5092		:	dataRd	 = 	 1'b0
;    5093		:	dataRd	 = 	 1'b0
;    5094		:	dataRd	 = 	 1'b0
;    5095		:	dataRd	 = 	 1'b0
;    5096		:	dataRd	 = 	 1'b0
;    5097		:	dataRd	 = 	 1'b0
;    5098		:	dataRd	 = 	 1'b0
;    5099		:	dataRd	 = 	 1'b0
;    5100		:	dataRd	 = 	 1'b0
;    5101		:	dataRd	 = 	 1'b0
;    5102		:	dataRd	 = 	 1'b0
;    5103		:	dataRd	 = 	 1'b0
;    5104		:	dataRd	 = 	 1'b0
;    5105		:	dataRd	 = 	 1'b0
;    5106		:	dataRd	 = 	 1'b0
;    5107		:	dataRd	 = 	 1'b0
;    5108		:	dataRd	 = 	 1'b0
;    5109		:	dataRd	 = 	 1'b0
;    5110		:	dataRd	 = 	 1'b0
;    5111		:	dataRd	 = 	 1'b0
;    5112		:	dataRd	 = 	 1'b0
;    5113		:	dataRd	 = 	 1'b0
;    5114		:	dataRd	 = 	 1'b0
;    5115		:	dataRd	 = 	 1'b0
;    5116		:	dataRd	 = 	 1'b0
;    5117		:	dataRd	 = 	 1'b0
;    5118		:	dataRd	 = 	 1'b0
;    5119		:	dataRd	 = 	 1'b0
;    5120		:	dataRd	 = 	 1'b0
;    5121		:	dataRd	 = 	 1'b0
;    5122		:	dataRd	 = 	 1'b0
;    5123		:	dataRd	 = 	 1'b0
;    5124		:	dataRd	 = 	 1'b0
;    5125		:	dataRd	 = 	 1'b0
;    5126		:	dataRd	 = 	 1'b0
;    5127		:	dataRd	 = 	 1'b0
;    5128		:	dataRd	 = 	 1'b0
;    5129		:	dataRd	 = 	 1'b0
;    5130		:	dataRd	 = 	 1'b0
;    5131		:	dataRd	 = 	 1'b0
;    5132		:	dataRd	 = 	 1'b0
;    5133		:	dataRd	 = 	 1'b0
;    5134		:	dataRd	 = 	 1'b0
;    5135		:	dataRd	 = 	 1'b0
;    5136		:	dataRd	 = 	 1'b0
;    5137		:	dataRd	 = 	 1'b0
;    5138		:	dataRd	 = 	 1'b0
;    5139		:	dataRd	 = 	 1'b0
;    5140		:	dataRd	 = 	 1'b0
;    5141		:	dataRd	 = 	 1'b0
;    5142		:	dataRd	 = 	 1'b0
;    5143		:	dataRd	 = 	 1'b0
;    5144		:	dataRd	 = 	 1'b0
;    5145		:	dataRd	 = 	 1'b0
;    5146		:	dataRd	 = 	 1'b0
;    5147		:	dataRd	 = 	 1'b0
;    5148		:	dataRd	 = 	 1'b0
;    5149		:	dataRd	 = 	 1'b0
;    5150		:	dataRd	 = 	 1'b0
;    5151		:	dataRd	 = 	 1'b0
;    5152		:	dataRd	 = 	 1'b0
;    5153		:	dataRd	 = 	 1'b0
;    5154		:	dataRd	 = 	 1'b1
;    5155		:	dataRd	 = 	 1'b1
;    5156		:	dataRd	 = 	 1'b0
;    5157		:	dataRd	 = 	 1'b0
;    5158		:	dataRd	 = 	 1'b0
;    5159		:	dataRd	 = 	 1'b0
;    5160		:	dataRd	 = 	 1'b0
;    5161		:	dataRd	 = 	 1'b0
;    5162		:	dataRd	 = 	 1'b0
;    5163		:	dataRd	 = 	 1'b0
;    5164		:	dataRd	 = 	 1'b1
;    5165		:	dataRd	 = 	 1'b0
;    5166		:	dataRd	 = 	 1'b0
;    5167		:	dataRd	 = 	 1'b0
;    5168		:	dataRd	 = 	 1'b1
;    5169		:	dataRd	 = 	 1'b1
;    5170		:	dataRd	 = 	 1'b0
;    5171		:	dataRd	 = 	 1'b0
;    5172		:	dataRd	 = 	 1'b0
;    5173		:	dataRd	 = 	 1'b0
;    5174		:	dataRd	 = 	 1'b0
;    5175		:	dataRd	 = 	 1'b1
;    5176		:	dataRd	 = 	 1'b0
;    5177		:	dataRd	 = 	 1'b0
;    5178		:	dataRd	 = 	 1'b0
;    5179		:	dataRd	 = 	 1'b0
;    5180		:	dataRd	 = 	 1'b0
;    5181		:	dataRd	 = 	 1'b0
;    5182		:	dataRd	 = 	 1'b0
;    5183		:	dataRd	 = 	 1'b0
;    5184		:	dataRd	 = 	 1'b0
;    5185		:	dataRd	 = 	 1'b0
;    5186		:	dataRd	 = 	 1'b0
;    5187		:	dataRd	 = 	 1'b0
;    5188		:	dataRd	 = 	 1'b1
;    5189		:	dataRd	 = 	 1'b1
;    5190		:	dataRd	 = 	 1'b0
;    5191		:	dataRd	 = 	 1'b0
;    5192		:	dataRd	 = 	 1'b1
;    5193		:	dataRd	 = 	 1'b0
;    5194		:	dataRd	 = 	 1'b0
;    5195		:	dataRd	 = 	 1'b0
;    5196		:	dataRd	 = 	 1'b0
;    5197		:	dataRd	 = 	 1'b0
;    5198		:	dataRd	 = 	 1'b1
;    5199		:	dataRd	 = 	 1'b0
;    5200		:	dataRd	 = 	 1'b0
;    5201		:	dataRd	 = 	 1'b0
;    5202		:	dataRd	 = 	 1'b0
;    5203		:	dataRd	 = 	 1'b0
;    5204		:	dataRd	 = 	 1'b0
;    5205		:	dataRd	 = 	 1'b0
;    5206		:	dataRd	 = 	 1'b0
;    5207		:	dataRd	 = 	 1'b0
;    5208		:	dataRd	 = 	 1'b0
;    5209		:	dataRd	 = 	 1'b0
;    5210		:	dataRd	 = 	 1'b0
;    5211		:	dataRd	 = 	 1'b0
;    5212		:	dataRd	 = 	 1'b0
;    5213		:	dataRd	 = 	 1'b0
;    5214		:	dataRd	 = 	 1'b1
;    5215		:	dataRd	 = 	 1'b0
;    5216		:	dataRd	 = 	 1'b0
;    5217		:	dataRd	 = 	 1'b0
;    5218		:	dataRd	 = 	 1'b0
;    5219		:	dataRd	 = 	 1'b0
;    5220		:	dataRd	 = 	 1'b0
;    5221		:	dataRd	 = 	 1'b0
;    5222		:	dataRd	 = 	 1'b0
;    5223		:	dataRd	 = 	 1'b0
;    5224		:	dataRd	 = 	 1'b0
;    5225		:	dataRd	 = 	 1'b0
;    5226		:	dataRd	 = 	 1'b0
;    5227		:	dataRd	 = 	 1'b0
;    5228		:	dataRd	 = 	 1'b0
;    5229		:	dataRd	 = 	 1'b0
;    5230		:	dataRd	 = 	 1'b1
;    5231		:	dataRd	 = 	 1'b0
;    5232		:	dataRd	 = 	 1'b0
;    5233		:	dataRd	 = 	 1'b0
;    5234		:	dataRd	 = 	 1'b0
;    5235		:	dataRd	 = 	 1'b0
;    5236		:	dataRd	 = 	 1'b0
;    5237		:	dataRd	 = 	 1'b0
;    5238		:	dataRd	 = 	 1'b0
;    5239		:	dataRd	 = 	 1'b0
;    5240		:	dataRd	 = 	 1'b0
;    5241		:	dataRd	 = 	 1'b0
;    5242		:	dataRd	 = 	 1'b0
;    5243		:	dataRd	 = 	 1'b0
;    5244		:	dataRd	 = 	 1'b0
;    5245		:	dataRd	 = 	 1'b0
;    5246		:	dataRd	 = 	 1'b1
;    5247		:	dataRd	 = 	 1'b0
;    5248		:	dataRd	 = 	 1'b0
;    5249		:	dataRd	 = 	 1'b0
;    5250		:	dataRd	 = 	 1'b0
;    5251		:	dataRd	 = 	 1'b0
;    5252		:	dataRd	 = 	 1'b0
;    5253		:	dataRd	 = 	 1'b0
;    5254		:	dataRd	 = 	 1'b0
;    5255		:	dataRd	 = 	 1'b0
;    5256		:	dataRd	 = 	 1'b0
;    5257		:	dataRd	 = 	 1'b0
;    5258		:	dataRd	 = 	 1'b0
;    5259		:	dataRd	 = 	 1'b0
;    5260		:	dataRd	 = 	 1'b0
;    5261		:	dataRd	 = 	 1'b0
;    5262		:	dataRd	 = 	 1'b1
;    5263		:	dataRd	 = 	 1'b0
;    5264		:	dataRd	 = 	 1'b0
;    5265		:	dataRd	 = 	 1'b0
;    5266		:	dataRd	 = 	 1'b0
;    5267		:	dataRd	 = 	 1'b0
;    5268		:	dataRd	 = 	 1'b0
;    5269		:	dataRd	 = 	 1'b0
;    5270		:	dataRd	 = 	 1'b0
;    5271		:	dataRd	 = 	 1'b0
;    5272		:	dataRd	 = 	 1'b0
;    5273		:	dataRd	 = 	 1'b0
;    5274		:	dataRd	 = 	 1'b0
;    5275		:	dataRd	 = 	 1'b0
;    5276		:	dataRd	 = 	 1'b0
;    5277		:	dataRd	 = 	 1'b0
;    5278		:	dataRd	 = 	 1'b1
;    5279		:	dataRd	 = 	 1'b0
;    5280		:	dataRd	 = 	 1'b0
;    5281		:	dataRd	 = 	 1'b0
;    5282		:	dataRd	 = 	 1'b0
;    5283		:	dataRd	 = 	 1'b0
;    5284		:	dataRd	 = 	 1'b0
;    5285		:	dataRd	 = 	 1'b0
;    5286		:	dataRd	 = 	 1'b0
;    5287		:	dataRd	 = 	 1'b0
;    5288		:	dataRd	 = 	 1'b0
;    5289		:	dataRd	 = 	 1'b0
;    5290		:	dataRd	 = 	 1'b0
;    5291		:	dataRd	 = 	 1'b0
;    5292		:	dataRd	 = 	 1'b0
;    5293		:	dataRd	 = 	 1'b0
;    5294		:	dataRd	 = 	 1'b1
;    5295		:	dataRd	 = 	 1'b0
;    5296		:	dataRd	 = 	 1'b0
;    5297		:	dataRd	 = 	 1'b0
;    5298		:	dataRd	 = 	 1'b0
;    5299		:	dataRd	 = 	 1'b0
;    5300		:	dataRd	 = 	 1'b0
;    5301		:	dataRd	 = 	 1'b0
;    5302		:	dataRd	 = 	 1'b0
;    5303		:	dataRd	 = 	 1'b0
;    5304		:	dataRd	 = 	 1'b0
;    5305		:	dataRd	 = 	 1'b0
;    5306		:	dataRd	 = 	 1'b0
;    5307		:	dataRd	 = 	 1'b0
;    5308		:	dataRd	 = 	 1'b0
;    5309		:	dataRd	 = 	 1'b0
;    5310		:	dataRd	 = 	 1'b1
;    5311		:	dataRd	 = 	 1'b0
;    5312		:	dataRd	 = 	 1'b0
;    5313		:	dataRd	 = 	 1'b0
;    5314		:	dataRd	 = 	 1'b0
;    5315		:	dataRd	 = 	 1'b0
;    5316		:	dataRd	 = 	 1'b0
;    5317		:	dataRd	 = 	 1'b0
;    5318		:	dataRd	 = 	 1'b0
;    5319		:	dataRd	 = 	 1'b0
;    5320		:	dataRd	 = 	 1'b0
;    5321		:	dataRd	 = 	 1'b0
;    5322		:	dataRd	 = 	 1'b0
;    5323		:	dataRd	 = 	 1'b0
;    5324		:	dataRd	 = 	 1'b0
;    5325		:	dataRd	 = 	 1'b0
;    5326		:	dataRd	 = 	 1'b1
;    5327		:	dataRd	 = 	 1'b0
;    5328		:	dataRd	 = 	 1'b0
;    5329		:	dataRd	 = 	 1'b0
;    5330		:	dataRd	 = 	 1'b0
;    5331		:	dataRd	 = 	 1'b0
;    5332		:	dataRd	 = 	 1'b0
;    5333		:	dataRd	 = 	 1'b0
;    5334		:	dataRd	 = 	 1'b0
;    5335		:	dataRd	 = 	 1'b0
;    5336		:	dataRd	 = 	 1'b0
;    5337		:	dataRd	 = 	 1'b0
;    5338		:	dataRd	 = 	 1'b0
;    5339		:	dataRd	 = 	 1'b0
;    5340		:	dataRd	 = 	 1'b0
;    5341		:	dataRd	 = 	 1'b0
;    5342		:	dataRd	 = 	 1'b1
;    5343		:	dataRd	 = 	 1'b0
;    5344		:	dataRd	 = 	 1'b0
;    5345		:	dataRd	 = 	 1'b0
;    5346		:	dataRd	 = 	 1'b0
;    5347		:	dataRd	 = 	 1'b0
;    5348		:	dataRd	 = 	 1'b0
;    5349		:	dataRd	 = 	 1'b0
;    5350		:	dataRd	 = 	 1'b0
;    5351		:	dataRd	 = 	 1'b0
;    5352		:	dataRd	 = 	 1'b0
;    5353		:	dataRd	 = 	 1'b0
;    5354		:	dataRd	 = 	 1'b0
;    5355		:	dataRd	 = 	 1'b0
;    5356		:	dataRd	 = 	 1'b0
;    5357		:	dataRd	 = 	 1'b0
;    5358		:	dataRd	 = 	 1'b1
;    5359		:	dataRd	 = 	 1'b0
;    5360		:	dataRd	 = 	 1'b0
;    5361		:	dataRd	 = 	 1'b0
;    5362		:	dataRd	 = 	 1'b0
;    5363		:	dataRd	 = 	 1'b0
;    5364		:	dataRd	 = 	 1'b0
;    5365		:	dataRd	 = 	 1'b0
;    5366		:	dataRd	 = 	 1'b0
;    5367		:	dataRd	 = 	 1'b0
;    5368		:	dataRd	 = 	 1'b0
;    5369		:	dataRd	 = 	 1'b0
;    5370		:	dataRd	 = 	 1'b0
;    5371		:	dataRd	 = 	 1'b0
;    5372		:	dataRd	 = 	 1'b0
;    5373		:	dataRd	 = 	 1'b0
;    5374		:	dataRd	 = 	 1'b1
;    5375		:	dataRd	 = 	 1'b0
;    5376		:	dataRd	 = 	 1'b0
;    5377		:	dataRd	 = 	 1'b0
;    5378		:	dataRd	 = 	 1'b0
;    5379		:	dataRd	 = 	 1'b0
;    5380		:	dataRd	 = 	 1'b0
;    5381		:	dataRd	 = 	 1'b0
;    5382		:	dataRd	 = 	 1'b0
;    5383		:	dataRd	 = 	 1'b0
;    5384		:	dataRd	 = 	 1'b0
;    5385		:	dataRd	 = 	 1'b0
;    5386		:	dataRd	 = 	 1'b0
;    5387		:	dataRd	 = 	 1'b0
;    5388		:	dataRd	 = 	 1'b0
;    5389		:	dataRd	 = 	 1'b0
;    5390		:	dataRd	 = 	 1'b1
;    5391		:	dataRd	 = 	 1'b0
;    5392		:	dataRd	 = 	 1'b0
;    5393		:	dataRd	 = 	 1'b0
;    5394		:	dataRd	 = 	 1'b0
;    5395		:	dataRd	 = 	 1'b0
;    5396		:	dataRd	 = 	 1'b0
;    5397		:	dataRd	 = 	 1'b0
;    5398		:	dataRd	 = 	 1'b0
;    5399		:	dataRd	 = 	 1'b0
;    5400		:	dataRd	 = 	 1'b0
;    5401		:	dataRd	 = 	 1'b0
;    5402		:	dataRd	 = 	 1'b0
;    5403		:	dataRd	 = 	 1'b0
;    5404		:	dataRd	 = 	 1'b0
;    5405		:	dataRd	 = 	 1'b0
;    5406		:	dataRd	 = 	 1'b1
;    5407		:	dataRd	 = 	 1'b0
;    5408		:	dataRd	 = 	 1'b0
;    5409		:	dataRd	 = 	 1'b0
;    5410		:	dataRd	 = 	 1'b0
;    5411		:	dataRd	 = 	 1'b0
;    5412		:	dataRd	 = 	 1'b0
;    5413		:	dataRd	 = 	 1'b0
;    5414		:	dataRd	 = 	 1'b0
;    5415		:	dataRd	 = 	 1'b0
;    5416		:	dataRd	 = 	 1'b0
;    5417		:	dataRd	 = 	 1'b0
;    5418		:	dataRd	 = 	 1'b0
;    5419		:	dataRd	 = 	 1'b0
;    5420		:	dataRd	 = 	 1'b0
;    5421		:	dataRd	 = 	 1'b0
;    5422		:	dataRd	 = 	 1'b1
;    5423		:	dataRd	 = 	 1'b0
;    5424		:	dataRd	 = 	 1'b0
;    5425		:	dataRd	 = 	 1'b0
;    5426		:	dataRd	 = 	 1'b0
;    5427		:	dataRd	 = 	 1'b0
;    5428		:	dataRd	 = 	 1'b0
;    5429		:	dataRd	 = 	 1'b0
;    5430		:	dataRd	 = 	 1'b0
;    5431		:	dataRd	 = 	 1'b0
;    5432		:	dataRd	 = 	 1'b0
;    5433		:	dataRd	 = 	 1'b0
;    5434		:	dataRd	 = 	 1'b0
;    5435		:	dataRd	 = 	 1'b0
;    5436		:	dataRd	 = 	 1'b0
;    5437		:	dataRd	 = 	 1'b0
;    5438		:	dataRd	 = 	 1'b1
;    5439		:	dataRd	 = 	 1'b0
;    5440		:	dataRd	 = 	 1'b0
;    5441		:	dataRd	 = 	 1'b0
;    5442		:	dataRd	 = 	 1'b0
;    5443		:	dataRd	 = 	 1'b0
;    5444		:	dataRd	 = 	 1'b0
;    5445		:	dataRd	 = 	 1'b0
;    5446		:	dataRd	 = 	 1'b0
;    5447		:	dataRd	 = 	 1'b0
;    5448		:	dataRd	 = 	 1'b0
;    5449		:	dataRd	 = 	 1'b0
;    5450		:	dataRd	 = 	 1'b0
;    5451		:	dataRd	 = 	 1'b0
;    5452		:	dataRd	 = 	 1'b0
;    5453		:	dataRd	 = 	 1'b0
;    5454		:	dataRd	 = 	 1'b1
;    5455		:	dataRd	 = 	 1'b0
;    5456		:	dataRd	 = 	 1'b0
;    5457		:	dataRd	 = 	 1'b0
;    5458		:	dataRd	 = 	 1'b0
;    5459		:	dataRd	 = 	 1'b0
;    5460		:	dataRd	 = 	 1'b0
;    5461		:	dataRd	 = 	 1'b0
;    5462		:	dataRd	 = 	 1'b0
;    5463		:	dataRd	 = 	 1'b0
;    5464		:	dataRd	 = 	 1'b0
;    5465		:	dataRd	 = 	 1'b0
;    5466		:	dataRd	 = 	 1'b0
;    5467		:	dataRd	 = 	 1'b0
;    5468		:	dataRd	 = 	 1'b0
;    5469		:	dataRd	 = 	 1'b0
;    5470		:	dataRd	 = 	 1'b1
;    5471		:	dataRd	 = 	 1'b0
;    5472		:	dataRd	 = 	 1'b0
;    5473		:	dataRd	 = 	 1'b0
;    5474		:	dataRd	 = 	 1'b0
;    5475		:	dataRd	 = 	 1'b0
;    5476		:	dataRd	 = 	 1'b0
;    5477		:	dataRd	 = 	 1'b0
;    5478		:	dataRd	 = 	 1'b0
;    5479		:	dataRd	 = 	 1'b0
;    5480		:	dataRd	 = 	 1'b0
;    5481		:	dataRd	 = 	 1'b0
;    5482		:	dataRd	 = 	 1'b0
;    5483		:	dataRd	 = 	 1'b0
;    5484		:	dataRd	 = 	 1'b0
;    5485		:	dataRd	 = 	 1'b0
;    5486		:	dataRd	 = 	 1'b1
;    5487		:	dataRd	 = 	 1'b0
;    5488		:	dataRd	 = 	 1'b0
;    5489		:	dataRd	 = 	 1'b0
;    5490		:	dataRd	 = 	 1'b0
;    5491		:	dataRd	 = 	 1'b0
;    5492		:	dataRd	 = 	 1'b0
;    5493		:	dataRd	 = 	 1'b0
;    5494		:	dataRd	 = 	 1'b0
;    5495		:	dataRd	 = 	 1'b0
;    5496		:	dataRd	 = 	 1'b0
;    5497		:	dataRd	 = 	 1'b0
;    5498		:	dataRd	 = 	 1'b0
;    5499		:	dataRd	 = 	 1'b0
;    5500		:	dataRd	 = 	 1'b0
;    5501		:	dataRd	 = 	 1'b0
;    5502		:	dataRd	 = 	 1'b1
;    5503		:	dataRd	 = 	 1'b0
;    5504		:	dataRd	 = 	 1'b0
;    5505		:	dataRd	 = 	 1'b0
;    5506		:	dataRd	 = 	 1'b0
;    5507		:	dataRd	 = 	 1'b0
;    5508		:	dataRd	 = 	 1'b0
;    5509		:	dataRd	 = 	 1'b0
;    5510		:	dataRd	 = 	 1'b0
;    5511		:	dataRd	 = 	 1'b0
;    5512		:	dataRd	 = 	 1'b0
;    5513		:	dataRd	 = 	 1'b0
;    5514		:	dataRd	 = 	 1'b0
;    5515		:	dataRd	 = 	 1'b0
;    5516		:	dataRd	 = 	 1'b0
;    5517		:	dataRd	 = 	 1'b0
;    5518		:	dataRd	 = 	 1'b1
;    5519		:	dataRd	 = 	 1'b0
;    5520		:	dataRd	 = 	 1'b0
;    5521		:	dataRd	 = 	 1'b0
;    5522		:	dataRd	 = 	 1'b0
;    5523		:	dataRd	 = 	 1'b0
;    5524		:	dataRd	 = 	 1'b0
;    5525		:	dataRd	 = 	 1'b0
;    5526		:	dataRd	 = 	 1'b0
;    5527		:	dataRd	 = 	 1'b0
;    5528		:	dataRd	 = 	 1'b0
;    5529		:	dataRd	 = 	 1'b0
;    5530		:	dataRd	 = 	 1'b0
;    5531		:	dataRd	 = 	 1'b0
;    5532		:	dataRd	 = 	 1'b0
;    5533		:	dataRd	 = 	 1'b0
;    5534		:	dataRd	 = 	 1'b1
;    5535		:	dataRd	 = 	 1'b0
;    5536		:	dataRd	 = 	 1'b0
;    5537		:	dataRd	 = 	 1'b0
;    5538		:	dataRd	 = 	 1'b0
;    5539		:	dataRd	 = 	 1'b0
;    5540		:	dataRd	 = 	 1'b0
;    5541		:	dataRd	 = 	 1'b0
;    5542		:	dataRd	 = 	 1'b0
;    5543		:	dataRd	 = 	 1'b0
;    5544		:	dataRd	 = 	 1'b0
;    5545		:	dataRd	 = 	 1'b0
;    5546		:	dataRd	 = 	 1'b0
;    5547		:	dataRd	 = 	 1'b0
;    5548		:	dataRd	 = 	 1'b0
;    5549		:	dataRd	 = 	 1'b0
;    5550		:	dataRd	 = 	 1'b1
;    5551		:	dataRd	 = 	 1'b0
;    5552		:	dataRd	 = 	 1'b0
;    5553		:	dataRd	 = 	 1'b0
;    5554		:	dataRd	 = 	 1'b0
;    5555		:	dataRd	 = 	 1'b0
;    5556		:	dataRd	 = 	 1'b0
;    5557		:	dataRd	 = 	 1'b0
;    5558		:	dataRd	 = 	 1'b0
;    5559		:	dataRd	 = 	 1'b0
;    5560		:	dataRd	 = 	 1'b0
;    5561		:	dataRd	 = 	 1'b0
;    5562		:	dataRd	 = 	 1'b0
;    5563		:	dataRd	 = 	 1'b0
;    5564		:	dataRd	 = 	 1'b0
;    5565		:	dataRd	 = 	 1'b0
;    5566		:	dataRd	 = 	 1'b1
;    5567		:	dataRd	 = 	 1'b0
;    5568		:	dataRd	 = 	 1'b0
;    5569		:	dataRd	 = 	 1'b0
;    5570		:	dataRd	 = 	 1'b0
;    5571		:	dataRd	 = 	 1'b0
;    5572		:	dataRd	 = 	 1'b0
;    5573		:	dataRd	 = 	 1'b0
;    5574		:	dataRd	 = 	 1'b0
;    5575		:	dataRd	 = 	 1'b0
;    5576		:	dataRd	 = 	 1'b0
;    5577		:	dataRd	 = 	 1'b0
;    5578		:	dataRd	 = 	 1'b0
;    5579		:	dataRd	 = 	 1'b0
;    5580		:	dataRd	 = 	 1'b0
;    5581		:	dataRd	 = 	 1'b0
;    5582		:	dataRd	 = 	 1'b1
;    5583		:	dataRd	 = 	 1'b0
;    5584		:	dataRd	 = 	 1'b0
;    5585		:	dataRd	 = 	 1'b0
;    5586		:	dataRd	 = 	 1'b0
;    5587		:	dataRd	 = 	 1'b0
;    5588		:	dataRd	 = 	 1'b0
;    5589		:	dataRd	 = 	 1'b0
;    5590		:	dataRd	 = 	 1'b0
;    5591		:	dataRd	 = 	 1'b0
;    5592		:	dataRd	 = 	 1'b0
;    5593		:	dataRd	 = 	 1'b0
;    5594		:	dataRd	 = 	 1'b0
;    5595		:	dataRd	 = 	 1'b0
;    5596		:	dataRd	 = 	 1'b0
;    5597		:	dataRd	 = 	 1'b0
;    5598		:	dataRd	 = 	 1'b1
;    5599		:	dataRd	 = 	 1'b0
;    5600		:	dataRd	 = 	 1'b0
;    5601		:	dataRd	 = 	 1'b0
;    5602		:	dataRd	 = 	 1'b0
;    5603		:	dataRd	 = 	 1'b0
;    5604		:	dataRd	 = 	 1'b0
;    5605		:	dataRd	 = 	 1'b0
;    5606		:	dataRd	 = 	 1'b0
;    5607		:	dataRd	 = 	 1'b0
;    5608		:	dataRd	 = 	 1'b0
;    5609		:	dataRd	 = 	 1'b0
;    5610		:	dataRd	 = 	 1'b0
;    5611		:	dataRd	 = 	 1'b0
;    5612		:	dataRd	 = 	 1'b0
;    5613		:	dataRd	 = 	 1'b0
;    5614		:	dataRd	 = 	 1'b1
;    5615		:	dataRd	 = 	 1'b0
;    5616		:	dataRd	 = 	 1'b0
;    5617		:	dataRd	 = 	 1'b0
;    5618		:	dataRd	 = 	 1'b0
;    5619		:	dataRd	 = 	 1'b0
;    5620		:	dataRd	 = 	 1'b0
;    5621		:	dataRd	 = 	 1'b0
;    5622		:	dataRd	 = 	 1'b0
;    5623		:	dataRd	 = 	 1'b0
;    5624		:	dataRd	 = 	 1'b0
;    5625		:	dataRd	 = 	 1'b0
;    5626		:	dataRd	 = 	 1'b0
;    5627		:	dataRd	 = 	 1'b0
;    5628		:	dataRd	 = 	 1'b0
;    5629		:	dataRd	 = 	 1'b0
;    5630		:	dataRd	 = 	 1'b1
;    5631		:	dataRd	 = 	 1'b0
;    5632		:	dataRd	 = 	 1'b0
;    5633		:	dataRd	 = 	 1'b0
;    5634		:	dataRd	 = 	 1'b0
;    5635		:	dataRd	 = 	 1'b0
;    5636		:	dataRd	 = 	 1'b0
;    5637		:	dataRd	 = 	 1'b0
;    5638		:	dataRd	 = 	 1'b0
;    5639		:	dataRd	 = 	 1'b0
;    5640		:	dataRd	 = 	 1'b0
;    5641		:	dataRd	 = 	 1'b0
;    5642		:	dataRd	 = 	 1'b0
;    5643		:	dataRd	 = 	 1'b0
;    5644		:	dataRd	 = 	 1'b0
;    5645		:	dataRd	 = 	 1'b0
;    5646		:	dataRd	 = 	 1'b1
;    5647		:	dataRd	 = 	 1'b0
;    5648		:	dataRd	 = 	 1'b0
;    5649		:	dataRd	 = 	 1'b0
;    5650		:	dataRd	 = 	 1'b0
;    5651		:	dataRd	 = 	 1'b0
;    5652		:	dataRd	 = 	 1'b0
;    5653		:	dataRd	 = 	 1'b0
;    5654		:	dataRd	 = 	 1'b0
;    5655		:	dataRd	 = 	 1'b0
;    5656		:	dataRd	 = 	 1'b0
;    5657		:	dataRd	 = 	 1'b0
;    5658		:	dataRd	 = 	 1'b0
;    5659		:	dataRd	 = 	 1'b0
;    5660		:	dataRd	 = 	 1'b0
;    5661		:	dataRd	 = 	 1'b0
;    5662		:	dataRd	 = 	 1'b1
;    5663		:	dataRd	 = 	 1'b0
;    5664		:	dataRd	 = 	 1'b0
;    5665		:	dataRd	 = 	 1'b0
;    5666		:	dataRd	 = 	 1'b0
;    5667		:	dataRd	 = 	 1'b0
;    5668		:	dataRd	 = 	 1'b0
;    5669		:	dataRd	 = 	 1'b0
;    5670		:	dataRd	 = 	 1'b0
;    5671		:	dataRd	 = 	 1'b0
;    5672		:	dataRd	 = 	 1'b0
;    5673		:	dataRd	 = 	 1'b0
;    5674		:	dataRd	 = 	 1'b0
;    5675		:	dataRd	 = 	 1'b0
;    5676		:	dataRd	 = 	 1'b0
;    5677		:	dataRd	 = 	 1'b0
;    5678		:	dataRd	 = 	 1'b1
;    5679		:	dataRd	 = 	 1'b0
;    5680		:	dataRd	 = 	 1'b0
;    5681		:	dataRd	 = 	 1'b0
;    5682		:	dataRd	 = 	 1'b0
;    5683		:	dataRd	 = 	 1'b0
;    5684		:	dataRd	 = 	 1'b0
;    5685		:	dataRd	 = 	 1'b0
;    5686		:	dataRd	 = 	 1'b0
;    5687		:	dataRd	 = 	 1'b0
;    5688		:	dataRd	 = 	 1'b0
;    5689		:	dataRd	 = 	 1'b0
;    5690		:	dataRd	 = 	 1'b0
;    5691		:	dataRd	 = 	 1'b0
;    5692		:	dataRd	 = 	 1'b0
;    5693		:	dataRd	 = 	 1'b0
;    5694		:	dataRd	 = 	 1'b1
;    5695		:	dataRd	 = 	 1'b0
;    5696		:	dataRd	 = 	 1'b0
;    5697		:	dataRd	 = 	 1'b0
;    5698		:	dataRd	 = 	 1'b0
;    5699		:	dataRd	 = 	 1'b0
;    5700		:	dataRd	 = 	 1'b0
;    5701		:	dataRd	 = 	 1'b0
;    5702		:	dataRd	 = 	 1'b0
;    5703		:	dataRd	 = 	 1'b0
;    5704		:	dataRd	 = 	 1'b0
;    5705		:	dataRd	 = 	 1'b0
;    5706		:	dataRd	 = 	 1'b0
;    5707		:	dataRd	 = 	 1'b0
;    5708		:	dataRd	 = 	 1'b0
;    5709		:	dataRd	 = 	 1'b0
;    5710		:	dataRd	 = 	 1'b1
;    5711		:	dataRd	 = 	 1'b0
;    5712		:	dataRd	 = 	 1'b0
;    5713		:	dataRd	 = 	 1'b0
;    5714		:	dataRd	 = 	 1'b0
;    5715		:	dataRd	 = 	 1'b0
;    5716		:	dataRd	 = 	 1'b0
;    5717		:	dataRd	 = 	 1'b0
;    5718		:	dataRd	 = 	 1'b0
;    5719		:	dataRd	 = 	 1'b0
;    5720		:	dataRd	 = 	 1'b0
;    5721		:	dataRd	 = 	 1'b0
;    5722		:	dataRd	 = 	 1'b0
;    5723		:	dataRd	 = 	 1'b0
;    5724		:	dataRd	 = 	 1'b0
;    5725		:	dataRd	 = 	 1'b0
;    5726		:	dataRd	 = 	 1'b1
;    5727		:	dataRd	 = 	 1'b0
;    5728		:	dataRd	 = 	 1'b0
;    5729		:	dataRd	 = 	 1'b0
;    5730		:	dataRd	 = 	 1'b0
;    5731		:	dataRd	 = 	 1'b0
;    5732		:	dataRd	 = 	 1'b0
;    5733		:	dataRd	 = 	 1'b0
;    5734		:	dataRd	 = 	 1'b0
;    5735		:	dataRd	 = 	 1'b0
;    5736		:	dataRd	 = 	 1'b0
;    5737		:	dataRd	 = 	 1'b0
;    5738		:	dataRd	 = 	 1'b0
;    5739		:	dataRd	 = 	 1'b0
;    5740		:	dataRd	 = 	 1'b0
;    5741		:	dataRd	 = 	 1'b0
;    5742		:	dataRd	 = 	 1'b1
;    5743		:	dataRd	 = 	 1'b0
;    5744		:	dataRd	 = 	 1'b0
;    5745		:	dataRd	 = 	 1'b0
;    5746		:	dataRd	 = 	 1'b0
;    5747		:	dataRd	 = 	 1'b0
;    5748		:	dataRd	 = 	 1'b0
;    5749		:	dataRd	 = 	 1'b0
;    5750		:	dataRd	 = 	 1'b0
;    5751		:	dataRd	 = 	 1'b0
;    5752		:	dataRd	 = 	 1'b0
;    5753		:	dataRd	 = 	 1'b0
;    5754		:	dataRd	 = 	 1'b0
;    5755		:	dataRd	 = 	 1'b0
;    5756		:	dataRd	 = 	 1'b0
;    5757		:	dataRd	 = 	 1'b0
;    5758		:	dataRd	 = 	 1'b1
;    5759		:	dataRd	 = 	 1'b0
;    5760		:	dataRd	 = 	 1'b0
;    5761		:	dataRd	 = 	 1'b0
;    5762		:	dataRd	 = 	 1'b0
;    5763		:	dataRd	 = 	 1'b0
;    5764		:	dataRd	 = 	 1'b0
;    5765		:	dataRd	 = 	 1'b0
;    5766		:	dataRd	 = 	 1'b0
;    5767		:	dataRd	 = 	 1'b0
;    5768		:	dataRd	 = 	 1'b0
;    5769		:	dataRd	 = 	 1'b0
;    5770		:	dataRd	 = 	 1'b0
;    5771		:	dataRd	 = 	 1'b0
;    5772		:	dataRd	 = 	 1'b0
;    5773		:	dataRd	 = 	 1'b0
;    5774		:	dataRd	 = 	 1'b1
;    5775		:	dataRd	 = 	 1'b0
;    5776		:	dataRd	 = 	 1'b0
;    5777		:	dataRd	 = 	 1'b0
;    5778		:	dataRd	 = 	 1'b0
;    5779		:	dataRd	 = 	 1'b0
;    5780		:	dataRd	 = 	 1'b0
;    5781		:	dataRd	 = 	 1'b0
;    5782		:	dataRd	 = 	 1'b0
;    5783		:	dataRd	 = 	 1'b0
;    5784		:	dataRd	 = 	 1'b0
;    5785		:	dataRd	 = 	 1'b0
;    5786		:	dataRd	 = 	 1'b0
;    5787		:	dataRd	 = 	 1'b0
;    5788		:	dataRd	 = 	 1'b0
;    5789		:	dataRd	 = 	 1'b0
;    5790		:	dataRd	 = 	 1'b1
;    5791		:	dataRd	 = 	 1'b0
;    5792		:	dataRd	 = 	 1'b0
;    5793		:	dataRd	 = 	 1'b0
;    5794		:	dataRd	 = 	 1'b0
;    5795		:	dataRd	 = 	 1'b0
;    5796		:	dataRd	 = 	 1'b0
;    5797		:	dataRd	 = 	 1'b0
;    5798		:	dataRd	 = 	 1'b0
;    5799		:	dataRd	 = 	 1'b0
;    5800		:	dataRd	 = 	 1'b0
;    5801		:	dataRd	 = 	 1'b0
;    5802		:	dataRd	 = 	 1'b0
;    5803		:	dataRd	 = 	 1'b0
;    5804		:	dataRd	 = 	 1'b0
;    5805		:	dataRd	 = 	 1'b0
;    5806		:	dataRd	 = 	 1'b1
;    5807		:	dataRd	 = 	 1'b0
;    5808		:	dataRd	 = 	 1'b0
;    5809		:	dataRd	 = 	 1'b0
;    5810		:	dataRd	 = 	 1'b0
;    5811		:	dataRd	 = 	 1'b0
;    5812		:	dataRd	 = 	 1'b0
;    5813		:	dataRd	 = 	 1'b0
;    5814		:	dataRd	 = 	 1'b0
;    5815		:	dataRd	 = 	 1'b0
;    5816		:	dataRd	 = 	 1'b0
;    5817		:	dataRd	 = 	 1'b0
;    5818		:	dataRd	 = 	 1'b0
;    5819		:	dataRd	 = 	 1'b0
;    5820		:	dataRd	 = 	 1'b0
;    5821		:	dataRd	 = 	 1'b0
;    5822		:	dataRd	 = 	 1'b1
;    5823		:	dataRd	 = 	 1'b0
;    5824		:	dataRd	 = 	 1'b0
;    5825		:	dataRd	 = 	 1'b0
;    5826		:	dataRd	 = 	 1'b0
;    5827		:	dataRd	 = 	 1'b0
;    5828		:	dataRd	 = 	 1'b0
;    5829		:	dataRd	 = 	 1'b0
;    5830		:	dataRd	 = 	 1'b0
;    5831		:	dataRd	 = 	 1'b0
;    5832		:	dataRd	 = 	 1'b0
;    5833		:	dataRd	 = 	 1'b0
;    5834		:	dataRd	 = 	 1'b0
;    5835		:	dataRd	 = 	 1'b0
;    5836		:	dataRd	 = 	 1'b0
;    5837		:	dataRd	 = 	 1'b0
;    5838		:	dataRd	 = 	 1'b1
;    5839		:	dataRd	 = 	 1'b0
;    5840		:	dataRd	 = 	 1'b0
;    5841		:	dataRd	 = 	 1'b0
;    5842		:	dataRd	 = 	 1'b0
;    5843		:	dataRd	 = 	 1'b0
;    5844		:	dataRd	 = 	 1'b0
;    5845		:	dataRd	 = 	 1'b0
;    5846		:	dataRd	 = 	 1'b0
;    5847		:	dataRd	 = 	 1'b0
;    5848		:	dataRd	 = 	 1'b0
;    5849		:	dataRd	 = 	 1'b0
;    5850		:	dataRd	 = 	 1'b0
;    5851		:	dataRd	 = 	 1'b0
;    5852		:	dataRd	 = 	 1'b0
;    5853		:	dataRd	 = 	 1'b0
;    5854		:	dataRd	 = 	 1'b1
;    5855		:	dataRd	 = 	 1'b0
;    5856		:	dataRd	 = 	 1'b0
;    5857		:	dataRd	 = 	 1'b0
;    5858		:	dataRd	 = 	 1'b0
;    5859		:	dataRd	 = 	 1'b0
;    5860		:	dataRd	 = 	 1'b0
;    5861		:	dataRd	 = 	 1'b0
;    5862		:	dataRd	 = 	 1'b0
;    5863		:	dataRd	 = 	 1'b0
;    5864		:	dataRd	 = 	 1'b0
;    5865		:	dataRd	 = 	 1'b0
;    5866		:	dataRd	 = 	 1'b0
;    5867		:	dataRd	 = 	 1'b0
;    5868		:	dataRd	 = 	 1'b0
;    5869		:	dataRd	 = 	 1'b0
;    5870		:	dataRd	 = 	 1'b1
;    5871		:	dataRd	 = 	 1'b0
;    5872		:	dataRd	 = 	 1'b0
;    5873		:	dataRd	 = 	 1'b0
;    5874		:	dataRd	 = 	 1'b0
;    5875		:	dataRd	 = 	 1'b0
;    5876		:	dataRd	 = 	 1'b0
;    5877		:	dataRd	 = 	 1'b0
;    5878		:	dataRd	 = 	 1'b0
;    5879		:	dataRd	 = 	 1'b0
;    5880		:	dataRd	 = 	 1'b0
;    5881		:	dataRd	 = 	 1'b0
;    5882		:	dataRd	 = 	 1'b0
;    5883		:	dataRd	 = 	 1'b0
;    5884		:	dataRd	 = 	 1'b0
;    5885		:	dataRd	 = 	 1'b0
;    5886		:	dataRd	 = 	 1'b1
;    5887		:	dataRd	 = 	 1'b0
;    5888		:	dataRd	 = 	 1'b0
;    5889		:	dataRd	 = 	 1'b0
;    5890		:	dataRd	 = 	 1'b0
;    5891		:	dataRd	 = 	 1'b0
;    5892		:	dataRd	 = 	 1'b0
;    5893		:	dataRd	 = 	 1'b0
;    5894		:	dataRd	 = 	 1'b0
;    5895		:	dataRd	 = 	 1'b0
;    5896		:	dataRd	 = 	 1'b0
;    5897		:	dataRd	 = 	 1'b0
;    5898		:	dataRd	 = 	 1'b0
;    5899		:	dataRd	 = 	 1'b0
;    5900		:	dataRd	 = 	 1'b0
;    5901		:	dataRd	 = 	 1'b0
;    5902		:	dataRd	 = 	 1'b1
;    5903		:	dataRd	 = 	 1'b0
;    5904		:	dataRd	 = 	 1'b0
;    5905		:	dataRd	 = 	 1'b0
;    5906		:	dataRd	 = 	 1'b0
;    5907		:	dataRd	 = 	 1'b0
;    5908		:	dataRd	 = 	 1'b0
;    5909		:	dataRd	 = 	 1'b0
;    5910		:	dataRd	 = 	 1'b0
;    5911		:	dataRd	 = 	 1'b0
;    5912		:	dataRd	 = 	 1'b0
;    5913		:	dataRd	 = 	 1'b0
;    5914		:	dataRd	 = 	 1'b0
;    5915		:	dataRd	 = 	 1'b0
;    5916		:	dataRd	 = 	 1'b0
;    5917		:	dataRd	 = 	 1'b0
;    5918		:	dataRd	 = 	 1'b1
;    5919		:	dataRd	 = 	 1'b0
;    5920		:	dataRd	 = 	 1'b0
;    5921		:	dataRd	 = 	 1'b0
;    5922		:	dataRd	 = 	 1'b0
;    5923		:	dataRd	 = 	 1'b0
;    5924		:	dataRd	 = 	 1'b0
;    5925		:	dataRd	 = 	 1'b0
;    5926		:	dataRd	 = 	 1'b0
;    5927		:	dataRd	 = 	 1'b0
;    5928		:	dataRd	 = 	 1'b0
;    5929		:	dataRd	 = 	 1'b0
;    5930		:	dataRd	 = 	 1'b0
;    5931		:	dataRd	 = 	 1'b0
;    5932		:	dataRd	 = 	 1'b0
;    5933		:	dataRd	 = 	 1'b0
;    5934		:	dataRd	 = 	 1'b1
;    5935		:	dataRd	 = 	 1'b0
;    5936		:	dataRd	 = 	 1'b0
;    5937		:	dataRd	 = 	 1'b0
;    5938		:	dataRd	 = 	 1'b0
;    5939		:	dataRd	 = 	 1'b0
;    5940		:	dataRd	 = 	 1'b0
;    5941		:	dataRd	 = 	 1'b0
;    5942		:	dataRd	 = 	 1'b0
;    5943		:	dataRd	 = 	 1'b0
;    5944		:	dataRd	 = 	 1'b0
;    5945		:	dataRd	 = 	 1'b0
;    5946		:	dataRd	 = 	 1'b0
;    5947		:	dataRd	 = 	 1'b0
;    5948		:	dataRd	 = 	 1'b0
;    5949		:	dataRd	 = 	 1'b0
;    5950		:	dataRd	 = 	 1'b1
;    5951		:	dataRd	 = 	 1'b0
;    5952		:	dataRd	 = 	 1'b0
;    5953		:	dataRd	 = 	 1'b0
;    5954		:	dataRd	 = 	 1'b0
;    5955		:	dataRd	 = 	 1'b0
;    5956		:	dataRd	 = 	 1'b0
;    5957		:	dataRd	 = 	 1'b0
;    5958		:	dataRd	 = 	 1'b0
;    5959		:	dataRd	 = 	 1'b0
;    5960		:	dataRd	 = 	 1'b0
;    5961		:	dataRd	 = 	 1'b0
;    5962		:	dataRd	 = 	 1'b0
;    5963		:	dataRd	 = 	 1'b0
;    5964		:	dataRd	 = 	 1'b0
;    5965		:	dataRd	 = 	 1'b0
;    5966		:	dataRd	 = 	 1'b1
;    5967		:	dataRd	 = 	 1'b0
;    5968		:	dataRd	 = 	 1'b0
;    5969		:	dataRd	 = 	 1'b0
;    5970		:	dataRd	 = 	 1'b0
;    5971		:	dataRd	 = 	 1'b0
;    5972		:	dataRd	 = 	 1'b0
;    5973		:	dataRd	 = 	 1'b0
;    5974		:	dataRd	 = 	 1'b0
;    5975		:	dataRd	 = 	 1'b0
;    5976		:	dataRd	 = 	 1'b0
;    5977		:	dataRd	 = 	 1'b0
;    5978		:	dataRd	 = 	 1'b0
;    5979		:	dataRd	 = 	 1'b0
;    5980		:	dataRd	 = 	 1'b0
;    5981		:	dataRd	 = 	 1'b0
;    5982		:	dataRd	 = 	 1'b1
;    5983		:	dataRd	 = 	 1'b0
;    5984		:	dataRd	 = 	 1'b0
;    5985		:	dataRd	 = 	 1'b0
;    5986		:	dataRd	 = 	 1'b0
;    5987		:	dataRd	 = 	 1'b0
;    5988		:	dataRd	 = 	 1'b0
;    5989		:	dataRd	 = 	 1'b0
;    5990		:	dataRd	 = 	 1'b0
;    5991		:	dataRd	 = 	 1'b0
;    5992		:	dataRd	 = 	 1'b0
;    5993		:	dataRd	 = 	 1'b0
;    5994		:	dataRd	 = 	 1'b0
;    5995		:	dataRd	 = 	 1'b0
;    5996		:	dataRd	 = 	 1'b0
;    5997		:	dataRd	 = 	 1'b0
;    5998		:	dataRd	 = 	 1'b1
;    5999		:	dataRd	 = 	 1'b0
;    6000		:	dataRd	 = 	 1'b0
;    6001		:	dataRd	 = 	 1'b0
;    6002		:	dataRd	 = 	 1'b0
;    6003		:	dataRd	 = 	 1'b0
;    6004		:	dataRd	 = 	 1'b0
;    6005		:	dataRd	 = 	 1'b0
;    6006		:	dataRd	 = 	 1'b0
;    6007		:	dataRd	 = 	 1'b0
;    6008		:	dataRd	 = 	 1'b0
;    6009		:	dataRd	 = 	 1'b0
;    6010		:	dataRd	 = 	 1'b0
;    6011		:	dataRd	 = 	 1'b0
;    6012		:	dataRd	 = 	 1'b0
;    6013		:	dataRd	 = 	 1'b0
;    6014		:	dataRd	 = 	 1'b1
;    6015		:	dataRd	 = 	 1'b0
;    6016		:	dataRd	 = 	 1'b0
;    6017		:	dataRd	 = 	 1'b0
;    6018		:	dataRd	 = 	 1'b0
;    6019		:	dataRd	 = 	 1'b0
;    6020		:	dataRd	 = 	 1'b0
;    6021		:	dataRd	 = 	 1'b0
;    6022		:	dataRd	 = 	 1'b0
;    6023		:	dataRd	 = 	 1'b0
;    6024		:	dataRd	 = 	 1'b0
;    6025		:	dataRd	 = 	 1'b0
;    6026		:	dataRd	 = 	 1'b0
;    6027		:	dataRd	 = 	 1'b0
;    6028		:	dataRd	 = 	 1'b0
;    6029		:	dataRd	 = 	 1'b0
;    6030		:	dataRd	 = 	 1'b1
;    6031		:	dataRd	 = 	 1'b0
;    6032		:	dataRd	 = 	 1'b0
;    6033		:	dataRd	 = 	 1'b0
;    6034		:	dataRd	 = 	 1'b0
;    6035		:	dataRd	 = 	 1'b0
;    6036		:	dataRd	 = 	 1'b0
;    6037		:	dataRd	 = 	 1'b0
;    6038		:	dataRd	 = 	 1'b0
;    6039		:	dataRd	 = 	 1'b0
;    6040		:	dataRd	 = 	 1'b0
;    6041		:	dataRd	 = 	 1'b0
;    6042		:	dataRd	 = 	 1'b0
;    6043		:	dataRd	 = 	 1'b0
;    6044		:	dataRd	 = 	 1'b0
;    6045		:	dataRd	 = 	 1'b0
;    6046		:	dataRd	 = 	 1'b1
;    6047		:	dataRd	 = 	 1'b0
;    6048		:	dataRd	 = 	 1'b0
;    6049		:	dataRd	 = 	 1'b0
;    6050		:	dataRd	 = 	 1'b0
;    6051		:	dataRd	 = 	 1'b0
;    6052		:	dataRd	 = 	 1'b0
;    6053		:	dataRd	 = 	 1'b0
;    6054		:	dataRd	 = 	 1'b0
;    6055		:	dataRd	 = 	 1'b0
;    6056		:	dataRd	 = 	 1'b0
;    6057		:	dataRd	 = 	 1'b0
;    6058		:	dataRd	 = 	 1'b0
;    6059		:	dataRd	 = 	 1'b0
;    6060		:	dataRd	 = 	 1'b0
;    6061		:	dataRd	 = 	 1'b0
;    6062		:	dataRd	 = 	 1'b1
;    6063		:	dataRd	 = 	 1'b0
;    6064		:	dataRd	 = 	 1'b0
;    6065		:	dataRd	 = 	 1'b0
;    6066		:	dataRd	 = 	 1'b0
;    6067		:	dataRd	 = 	 1'b0
;    6068		:	dataRd	 = 	 1'b0
;    6069		:	dataRd	 = 	 1'b0
;    6070		:	dataRd	 = 	 1'b0
;    6071		:	dataRd	 = 	 1'b0
;    6072		:	dataRd	 = 	 1'b0
;    6073		:	dataRd	 = 	 1'b0
;    6074		:	dataRd	 = 	 1'b0
;    6075		:	dataRd	 = 	 1'b0
;    6076		:	dataRd	 = 	 1'b0
;    6077		:	dataRd	 = 	 1'b0
;    6078		:	dataRd	 = 	 1'b1
;    6079		:	dataRd	 = 	 1'b0
;    6080		:	dataRd	 = 	 1'b0
;    6081		:	dataRd	 = 	 1'b0
;    6082		:	dataRd	 = 	 1'b0
;    6083		:	dataRd	 = 	 1'b0
;    6084		:	dataRd	 = 	 1'b0
;    6085		:	dataRd	 = 	 1'b0
;    6086		:	dataRd	 = 	 1'b0
;    6087		:	dataRd	 = 	 1'b0
;    6088		:	dataRd	 = 	 1'b0
;    6089		:	dataRd	 = 	 1'b0
;    6090		:	dataRd	 = 	 1'b0
;    6091		:	dataRd	 = 	 1'b0
;    6092		:	dataRd	 = 	 1'b0
;    6093		:	dataRd	 = 	 1'b0
;    6094		:	dataRd	 = 	 1'b1
;    6095		:	dataRd	 = 	 1'b0
;    6096		:	dataRd	 = 	 1'b0
;    6097		:	dataRd	 = 	 1'b0
;    6098		:	dataRd	 = 	 1'b0
;    6099		:	dataRd	 = 	 1'b0
;    6100		:	dataRd	 = 	 1'b0
;    6101		:	dataRd	 = 	 1'b0
;    6102		:	dataRd	 = 	 1'b0
;    6103		:	dataRd	 = 	 1'b0
;    6104		:	dataRd	 = 	 1'b0
;    6105		:	dataRd	 = 	 1'b0
;    6106		:	dataRd	 = 	 1'b0
;    6107		:	dataRd	 = 	 1'b0
;    6108		:	dataRd	 = 	 1'b0
;    6109		:	dataRd	 = 	 1'b0
;    6110		:	dataRd	 = 	 1'b1
;    6111		:	dataRd	 = 	 1'b0
;    6112		:	dataRd	 = 	 1'b0
;    6113		:	dataRd	 = 	 1'b0
;    6114		:	dataRd	 = 	 1'b0
;    6115		:	dataRd	 = 	 1'b0
;    6116		:	dataRd	 = 	 1'b0
;    6117		:	dataRd	 = 	 1'b0
;    6118		:	dataRd	 = 	 1'b0
;    6119		:	dataRd	 = 	 1'b0
;    6120		:	dataRd	 = 	 1'b0
;    6121		:	dataRd	 = 	 1'b0
;    6122		:	dataRd	 = 	 1'b0
;    6123		:	dataRd	 = 	 1'b0
;    6124		:	dataRd	 = 	 1'b0
;    6125		:	dataRd	 = 	 1'b0
;    6126		:	dataRd	 = 	 1'b1
;    6127		:	dataRd	 = 	 1'b0
;    6128		:	dataRd	 = 	 1'b0
;    6129		:	dataRd	 = 	 1'b0
;    6130		:	dataRd	 = 	 1'b0
;    6131		:	dataRd	 = 	 1'b0
;    6132		:	dataRd	 = 	 1'b0
;    6133		:	dataRd	 = 	 1'b0
;    6134		:	dataRd	 = 	 1'b0
;    6135		:	dataRd	 = 	 1'b0
;    6136		:	dataRd	 = 	 1'b0
;    6137		:	dataRd	 = 	 1'b0
;    6138		:	dataRd	 = 	 1'b0
;    6139		:	dataRd	 = 	 1'b0
;    6140		:	dataRd	 = 	 1'b0
;    6141		:	dataRd	 = 	 1'b0
;    6142		:	dataRd	 = 	 1'b1
;    6143		:	dataRd	 = 	 1'b0
;    6144		:	dataRd	 = 	 1'b0
;    6145		:	dataRd	 = 	 1'b0
;    6146		:	dataRd	 = 	 1'b0
;    6147		:	dataRd	 = 	 1'b0
;    6148		:	dataRd	 = 	 1'b0
;    6149		:	dataRd	 = 	 1'b0
;    6150		:	dataRd	 = 	 1'b0
;    6151		:	dataRd	 = 	 1'b0
;    6152		:	dataRd	 = 	 1'b0
;    6153		:	dataRd	 = 	 1'b0
;    6154		:	dataRd	 = 	 1'b0
;    6155		:	dataRd	 = 	 1'b0
;    6156		:	dataRd	 = 	 1'b0
;    6157		:	dataRd	 = 	 1'b0
;    6158		:	dataRd	 = 	 1'b1
;    6159		:	dataRd	 = 	 1'b0
;    6160		:	dataRd	 = 	 1'b0
;    6161		:	dataRd	 = 	 1'b0
;    6162		:	dataRd	 = 	 1'b0
;    6163		:	dataRd	 = 	 1'b0
;    6164		:	dataRd	 = 	 1'b0
;    6165		:	dataRd	 = 	 1'b0
;    6166		:	dataRd	 = 	 1'b0
;    6167		:	dataRd	 = 	 1'b0
;    6168		:	dataRd	 = 	 1'b0
;    6169		:	dataRd	 = 	 1'b0
;    6170		:	dataRd	 = 	 1'b0
;    6171		:	dataRd	 = 	 1'b0
;    6172		:	dataRd	 = 	 1'b0
;    6173		:	dataRd	 = 	 1'b0
;    6174		:	dataRd	 = 	 1'b0
;    6175		:	dataRd	 = 	 1'b0
;    6176		:	dataRd	 = 	 1'b0
;    6177		:	dataRd	 = 	 1'b0
;    6178		:	dataRd	 = 	 1'b0
;    6179		:	dataRd	 = 	 1'b0
;    6180		:	dataRd	 = 	 1'b0
;    6181		:	dataRd	 = 	 1'b0
;    6182		:	dataRd	 = 	 1'b0
;    6183		:	dataRd	 = 	 1'b0
;    6184		:	dataRd	 = 	 1'b0
;    6185		:	dataRd	 = 	 1'b0
;    6186		:	dataRd	 = 	 1'b0
;    6187		:	dataRd	 = 	 1'b0
;    6188		:	dataRd	 = 	 1'b0
;    6189		:	dataRd	 = 	 1'b0
;    6190		:	dataRd	 = 	 1'b0
;    6191		:	dataRd	 = 	 1'b0
;    6192		:	dataRd	 = 	 1'b0
;    6193		:	dataRd	 = 	 1'b0
;    6194		:	dataRd	 = 	 1'b0
;    6195		:	dataRd	 = 	 1'b0
;    6196		:	dataRd	 = 	 1'b0
;    6197		:	dataRd	 = 	 1'b0
;    6198		:	dataRd	 = 	 1'b0
;    6199		:	dataRd	 = 	 1'b0
;    6200		:	dataRd	 = 	 1'b0
;    6201		:	dataRd	 = 	 1'b0
;    6202		:	dataRd	 = 	 1'b0
;    6203		:	dataRd	 = 	 1'b0
;    6204		:	dataRd	 = 	 1'b0
;    6205		:	dataRd	 = 	 1'b0
;    6206		:	dataRd	 = 	 1'b0
;    6207		:	dataRd	 = 	 1'b0
;    6208		:	dataRd	 = 	 1'b0
;    6209		:	dataRd	 = 	 1'b0
;    6210		:	dataRd	 = 	 1'b0
;    6211		:	dataRd	 = 	 1'b0
;    6212		:	dataRd	 = 	 1'b0
;    6213		:	dataRd	 = 	 1'b0
;    6214		:	dataRd	 = 	 1'b0
;    6215		:	dataRd	 = 	 1'b0
;    6216		:	dataRd	 = 	 1'b0
;    6217		:	dataRd	 = 	 1'b0
;    6218		:	dataRd	 = 	 1'b0
;    6219		:	dataRd	 = 	 1'b0
;    6220		:	dataRd	 = 	 1'b0
;    6221		:	dataRd	 = 	 1'b0
;    6222		:	dataRd	 = 	 1'b0
;    6223		:	dataRd	 = 	 1'b0
;    6224		:	dataRd	 = 	 1'b0
;    6225		:	dataRd	 = 	 1'b1
;    6226		:	dataRd	 = 	 1'b0
;    6227		:	dataRd	 = 	 1'b0
;    6228		:	dataRd	 = 	 1'b0
;    6229		:	dataRd	 = 	 1'b0
;    6230		:	dataRd	 = 	 1'b0
;    6231		:	dataRd	 = 	 1'b0
;    6232		:	dataRd	 = 	 1'b0
;    6233		:	dataRd	 = 	 1'b0
;    6234		:	dataRd	 = 	 1'b0
;    6235		:	dataRd	 = 	 1'b0
;    6236		:	dataRd	 = 	 1'b0
;    6237		:	dataRd	 = 	 1'b0
;    6238		:	dataRd	 = 	 1'b0
;    6239		:	dataRd	 = 	 1'b0
;    6240		:	dataRd	 = 	 1'b0
;    6241		:	dataRd	 = 	 1'b0
;    6242		:	dataRd	 = 	 1'b0
;    6243		:	dataRd	 = 	 1'b0
;    6244		:	dataRd	 = 	 1'b0
;    6245		:	dataRd	 = 	 1'b0
;    6246		:	dataRd	 = 	 1'b0
;    6247		:	dataRd	 = 	 1'b0
;    6248		:	dataRd	 = 	 1'b0
;    6249		:	dataRd	 = 	 1'b0
;    6250		:	dataRd	 = 	 1'b0
;    6251		:	dataRd	 = 	 1'b0
;    6252		:	dataRd	 = 	 1'b0
;    6253		:	dataRd	 = 	 1'b0
;    6254		:	dataRd	 = 	 1'b0
;    6255		:	dataRd	 = 	 1'b0
;    6256		:	dataRd	 = 	 1'b0
;    6257		:	dataRd	 = 	 1'b0
;    6258		:	dataRd	 = 	 1'b0
;    6259		:	dataRd	 = 	 1'b0
;    6260		:	dataRd	 = 	 1'b0
;    6261		:	dataRd	 = 	 1'b0
;    6262		:	dataRd	 = 	 1'b0
;    6263		:	dataRd	 = 	 1'b0
;    6264		:	dataRd	 = 	 1'b0
;    6265		:	dataRd	 = 	 1'b0
;    6266		:	dataRd	 = 	 1'b0
;    6267		:	dataRd	 = 	 1'b0
;    6268		:	dataRd	 = 	 1'b0
;    6269		:	dataRd	 = 	 1'b0
;    6270		:	dataRd	 = 	 1'b0
;    6271		:	dataRd	 = 	 1'b0
;    6272		:	dataRd	 = 	 1'b0
;    6273		:	dataRd	 = 	 1'b0
;    6274		:	dataRd	 = 	 1'b0
;    6275		:	dataRd	 = 	 1'b0
;    6276		:	dataRd	 = 	 1'b0
;    6277		:	dataRd	 = 	 1'b0
;    6278		:	dataRd	 = 	 1'b0
;    6279		:	dataRd	 = 	 1'b0
;    6280		:	dataRd	 = 	 1'b0
;    6281		:	dataRd	 = 	 1'b0
;    6282		:	dataRd	 = 	 1'b0
;    6283		:	dataRd	 = 	 1'b0
;    6284		:	dataRd	 = 	 1'b0
;    6285		:	dataRd	 = 	 1'b0
;    6286		:	dataRd	 = 	 1'b0
;    6287		:	dataRd	 = 	 1'b0
;    6288		:	dataRd	 = 	 1'b0
;    6289		:	dataRd	 = 	 1'b0
;    6290		:	dataRd	 = 	 1'b0
;    6291		:	dataRd	 = 	 1'b0
;    6292		:	dataRd	 = 	 1'b1
;    6293		:	dataRd	 = 	 1'b0
;    6294		:	dataRd	 = 	 1'b0
;    6295		:	dataRd	 = 	 1'b0
;    6296		:	dataRd	 = 	 1'b0
;    6297		:	dataRd	 = 	 1'b0
;    6298		:	dataRd	 = 	 1'b0
;    6299		:	dataRd	 = 	 1'b0
;    6300		:	dataRd	 = 	 1'b0
;    6301		:	dataRd	 = 	 1'b0
;    6302		:	dataRd	 = 	 1'b0
;    6303		:	dataRd	 = 	 1'b0
;    6304		:	dataRd	 = 	 1'b0
;    6305		:	dataRd	 = 	 1'b0
;    6306		:	dataRd	 = 	 1'b0
;    6307		:	dataRd	 = 	 1'b0
;    6308		:	dataRd	 = 	 1'b0
;    6309		:	dataRd	 = 	 1'b0
;    6310		:	dataRd	 = 	 1'b0
;    6311		:	dataRd	 = 	 1'b0
;    6312		:	dataRd	 = 	 1'b0
;    6313		:	dataRd	 = 	 1'b0
;    6314		:	dataRd	 = 	 1'b0
;    6315		:	dataRd	 = 	 1'b0
;    6316		:	dataRd	 = 	 1'b0
;    6317		:	dataRd	 = 	 1'b0
;    6318		:	dataRd	 = 	 1'b0
;    6319		:	dataRd	 = 	 1'b0
;    6320		:	dataRd	 = 	 1'b0
;    6321		:	dataRd	 = 	 1'b0
;    6322		:	dataRd	 = 	 1'b0
;    6323		:	dataRd	 = 	 1'b0
;    6324		:	dataRd	 = 	 1'b0
;    6325		:	dataRd	 = 	 1'b0
;    6326		:	dataRd	 = 	 1'b0
;    6327		:	dataRd	 = 	 1'b0
;    6328		:	dataRd	 = 	 1'b0
;    6329		:	dataRd	 = 	 1'b0
;    6330		:	dataRd	 = 	 1'b0
;    6331		:	dataRd	 = 	 1'b0
;    6332		:	dataRd	 = 	 1'b0
;    6333		:	dataRd	 = 	 1'b0
;    6334		:	dataRd	 = 	 1'b0
;    6335		:	dataRd	 = 	 1'b0
;    6336		:	dataRd	 = 	 1'b0
;    6337		:	dataRd	 = 	 1'b0
;    6338		:	dataRd	 = 	 1'b0
;    6339		:	dataRd	 = 	 1'b0
;    6340		:	dataRd	 = 	 1'b0
;    6341		:	dataRd	 = 	 1'b0
;    6342		:	dataRd	 = 	 1'b0
;    6343		:	dataRd	 = 	 1'b0
;    6344		:	dataRd	 = 	 1'b0
;    6345		:	dataRd	 = 	 1'b0
;    6346		:	dataRd	 = 	 1'b0
;    6347		:	dataRd	 = 	 1'b0
;    6348		:	dataRd	 = 	 1'b0
;    6349		:	dataRd	 = 	 1'b0
;    6350		:	dataRd	 = 	 1'b0
;    6351		:	dataRd	 = 	 1'b0
;    6352		:	dataRd	 = 	 1'b0
;    6353		:	dataRd	 = 	 1'b0
;    6354		:	dataRd	 = 	 1'b0
;    6355		:	dataRd	 = 	 1'b0
;    6356		:	dataRd	 = 	 1'b0
;    6357		:	dataRd	 = 	 1'b0
;    6358		:	dataRd	 = 	 1'b0
;    6359		:	dataRd	 = 	 1'b1
;    6360		:	dataRd	 = 	 1'b0
;    6361		:	dataRd	 = 	 1'b0
;    6362		:	dataRd	 = 	 1'b0
;    6363		:	dataRd	 = 	 1'b0
;    6364		:	dataRd	 = 	 1'b0
;    6365		:	dataRd	 = 	 1'b0
;    6366		:	dataRd	 = 	 1'b0
;    6367		:	dataRd	 = 	 1'b0
;    6368		:	dataRd	 = 	 1'b0
;    6369		:	dataRd	 = 	 1'b0
;    6370		:	dataRd	 = 	 1'b0
;    6371		:	dataRd	 = 	 1'b0
;    6372		:	dataRd	 = 	 1'b0
;    6373		:	dataRd	 = 	 1'b0
;    6374		:	dataRd	 = 	 1'b0
;    6375		:	dataRd	 = 	 1'b0
;    6376		:	dataRd	 = 	 1'b0
;    6377		:	dataRd	 = 	 1'b0
;    6378		:	dataRd	 = 	 1'b0
;    6379		:	dataRd	 = 	 1'b0
;    6380		:	dataRd	 = 	 1'b0
;    6381		:	dataRd	 = 	 1'b0
;    6382		:	dataRd	 = 	 1'b0
;    6383		:	dataRd	 = 	 1'b0
;    6384		:	dataRd	 = 	 1'b0
;    6385		:	dataRd	 = 	 1'b0
;    6386		:	dataRd	 = 	 1'b0
;    6387		:	dataRd	 = 	 1'b0
;    6388		:	dataRd	 = 	 1'b0
;    6389		:	dataRd	 = 	 1'b0
;    6390		:	dataRd	 = 	 1'b0
;    6391		:	dataRd	 = 	 1'b0
;    6392		:	dataRd	 = 	 1'b0
;    6393		:	dataRd	 = 	 1'b0
;    6394		:	dataRd	 = 	 1'b0
;    6395		:	dataRd	 = 	 1'b0
;    6396		:	dataRd	 = 	 1'b0
;    6397		:	dataRd	 = 	 1'b0
;    6398		:	dataRd	 = 	 1'b0
;    6399		:	dataRd	 = 	 1'b0
;    6400		:	dataRd	 = 	 1'b0
;    6401		:	dataRd	 = 	 1'b0
;    6402		:	dataRd	 = 	 1'b0
;    6403		:	dataRd	 = 	 1'b0
;    6404		:	dataRd	 = 	 1'b0
;    6405		:	dataRd	 = 	 1'b0
;    6406		:	dataRd	 = 	 1'b0
;    6407		:	dataRd	 = 	 1'b0
;    6408		:	dataRd	 = 	 1'b0
;    6409		:	dataRd	 = 	 1'b0
;    6410		:	dataRd	 = 	 1'b0
;    6411		:	dataRd	 = 	 1'b0
;    6412		:	dataRd	 = 	 1'b0
;    6413		:	dataRd	 = 	 1'b0
;    6414		:	dataRd	 = 	 1'b0
;    6415		:	dataRd	 = 	 1'b0
;    6416		:	dataRd	 = 	 1'b0
;    6417		:	dataRd	 = 	 1'b0
;    6418		:	dataRd	 = 	 1'b0
;    6419		:	dataRd	 = 	 1'b0
;    6420		:	dataRd	 = 	 1'b0
;    6421		:	dataRd	 = 	 1'b0
;    6422		:	dataRd	 = 	 1'b0
;    6423		:	dataRd	 = 	 1'b0
;    6424		:	dataRd	 = 	 1'b0
;    6425		:	dataRd	 = 	 1'b0
;    6426		:	dataRd	 = 	 1'b1
;    6427		:	dataRd	 = 	 1'b0
;    6428		:	dataRd	 = 	 1'b0
;    6429		:	dataRd	 = 	 1'b0
;    6430		:	dataRd	 = 	 1'b0
;    6431		:	dataRd	 = 	 1'b0
;    6432		:	dataRd	 = 	 1'b0
;    6433		:	dataRd	 = 	 1'b0
;    6434		:	dataRd	 = 	 1'b0
;    6435		:	dataRd	 = 	 1'b0
;    6436		:	dataRd	 = 	 1'b0
;    6437		:	dataRd	 = 	 1'b0
;    6438		:	dataRd	 = 	 1'b0
;    6439		:	dataRd	 = 	 1'b0
;    6440		:	dataRd	 = 	 1'b0
;    6441		:	dataRd	 = 	 1'b0
;    6442		:	dataRd	 = 	 1'b0
;    6443		:	dataRd	 = 	 1'b0
;    6444		:	dataRd	 = 	 1'b0
;    6445		:	dataRd	 = 	 1'b0
;    6446		:	dataRd	 = 	 1'b0
;    6447		:	dataRd	 = 	 1'b0
;    6448		:	dataRd	 = 	 1'b0
;    6449		:	dataRd	 = 	 1'b0
;    6450		:	dataRd	 = 	 1'b0
;    6451		:	dataRd	 = 	 1'b0
;    6452		:	dataRd	 = 	 1'b0
;    6453		:	dataRd	 = 	 1'b0
;    6454		:	dataRd	 = 	 1'b0
;    6455		:	dataRd	 = 	 1'b0
;    6456		:	dataRd	 = 	 1'b0
;    6457		:	dataRd	 = 	 1'b0
;    6458		:	dataRd	 = 	 1'b0
;    6459		:	dataRd	 = 	 1'b0
;    6460		:	dataRd	 = 	 1'b0
;    6461		:	dataRd	 = 	 1'b0
;    6462		:	dataRd	 = 	 1'b0
;    6463		:	dataRd	 = 	 1'b0
;    6464		:	dataRd	 = 	 1'b0
;    6465		:	dataRd	 = 	 1'b0
;    6466		:	dataRd	 = 	 1'b0
;    6467		:	dataRd	 = 	 1'b0
;    6468		:	dataRd	 = 	 1'b0
;    6469		:	dataRd	 = 	 1'b0
;    6470		:	dataRd	 = 	 1'b0
;    6471		:	dataRd	 = 	 1'b0
;    6472		:	dataRd	 = 	 1'b0
;    6473		:	dataRd	 = 	 1'b0
;    6474		:	dataRd	 = 	 1'b0
;    6475		:	dataRd	 = 	 1'b0
;    6476		:	dataRd	 = 	 1'b0
;    6477		:	dataRd	 = 	 1'b0
;    6478		:	dataRd	 = 	 1'b0
;    6479		:	dataRd	 = 	 1'b0
;    6480		:	dataRd	 = 	 1'b0
;    6481		:	dataRd	 = 	 1'b0
;    6482		:	dataRd	 = 	 1'b0
;    6483		:	dataRd	 = 	 1'b0
;    6484		:	dataRd	 = 	 1'b0
;    6485		:	dataRd	 = 	 1'b0
;    6486		:	dataRd	 = 	 1'b0
;    6487		:	dataRd	 = 	 1'b0
;    6488		:	dataRd	 = 	 1'b0
;    6489		:	dataRd	 = 	 1'b0
;    6490		:	dataRd	 = 	 1'b0
;    6491		:	dataRd	 = 	 1'b0
;    6492		:	dataRd	 = 	 1'b0
;    6493		:	dataRd	 = 	 1'b1
;    6494		:	dataRd	 = 	 1'b0
;    6495		:	dataRd	 = 	 1'b0
;    6496		:	dataRd	 = 	 1'b0
;    6497		:	dataRd	 = 	 1'b0
;    6498		:	dataRd	 = 	 1'b0
;    6499		:	dataRd	 = 	 1'b0
;    6500		:	dataRd	 = 	 1'b0
;    6501		:	dataRd	 = 	 1'b0
;    6502		:	dataRd	 = 	 1'b0
;    6503		:	dataRd	 = 	 1'b0
;    6504		:	dataRd	 = 	 1'b0
;    6505		:	dataRd	 = 	 1'b0
;    6506		:	dataRd	 = 	 1'b0
;    6507		:	dataRd	 = 	 1'b0
;    6508		:	dataRd	 = 	 1'b0
;    6509		:	dataRd	 = 	 1'b0
;    6510		:	dataRd	 = 	 1'b0
;    6511		:	dataRd	 = 	 1'b0
;    6512		:	dataRd	 = 	 1'b0
;    6513		:	dataRd	 = 	 1'b0
;    6514		:	dataRd	 = 	 1'b0
;    6515		:	dataRd	 = 	 1'b0
;    6516		:	dataRd	 = 	 1'b0
;    6517		:	dataRd	 = 	 1'b0
;    6518		:	dataRd	 = 	 1'b0
;    6519		:	dataRd	 = 	 1'b0
;    6520		:	dataRd	 = 	 1'b0
;    6521		:	dataRd	 = 	 1'b0
;    6522		:	dataRd	 = 	 1'b0
;    6523		:	dataRd	 = 	 1'b0
;    6524		:	dataRd	 = 	 1'b0
;    6525		:	dataRd	 = 	 1'b0
;    6526		:	dataRd	 = 	 1'b0
;    6527		:	dataRd	 = 	 1'b0
;    6528		:	dataRd	 = 	 1'b0
;    6529		:	dataRd	 = 	 1'b0
;    6530		:	dataRd	 = 	 1'b0
;    6531		:	dataRd	 = 	 1'b0
;    6532		:	dataRd	 = 	 1'b0
;    6533		:	dataRd	 = 	 1'b0
;    6534		:	dataRd	 = 	 1'b0
;    6535		:	dataRd	 = 	 1'b0
;    6536		:	dataRd	 = 	 1'b0
;    6537		:	dataRd	 = 	 1'b0
;    6538		:	dataRd	 = 	 1'b0
;    6539		:	dataRd	 = 	 1'b0
;    6540		:	dataRd	 = 	 1'b0
;    6541		:	dataRd	 = 	 1'b0
;    6542		:	dataRd	 = 	 1'b0
;    6543		:	dataRd	 = 	 1'b0
;    6544		:	dataRd	 = 	 1'b0
;    6545		:	dataRd	 = 	 1'b0
;    6546		:	dataRd	 = 	 1'b0
;    6547		:	dataRd	 = 	 1'b0
;    6548		:	dataRd	 = 	 1'b0
;    6549		:	dataRd	 = 	 1'b0
;    6550		:	dataRd	 = 	 1'b0
;    6551		:	dataRd	 = 	 1'b0
;    6552		:	dataRd	 = 	 1'b0
;    6553		:	dataRd	 = 	 1'b0
;    6554		:	dataRd	 = 	 1'b0
;    6555		:	dataRd	 = 	 1'b0
;    6556		:	dataRd	 = 	 1'b0
;    6557		:	dataRd	 = 	 1'b0
;    6558		:	dataRd	 = 	 1'b0
;    6559		:	dataRd	 = 	 1'b0
;    6560		:	dataRd	 = 	 1'b1
;    6561		:	dataRd	 = 	 1'b0
;    6562		:	dataRd	 = 	 1'b0
;    6563		:	dataRd	 = 	 1'b0
;    6564		:	dataRd	 = 	 1'b0
;    6565		:	dataRd	 = 	 1'b0
;    6566		:	dataRd	 = 	 1'b0
;    6567		:	dataRd	 = 	 1'b0
;    6568		:	dataRd	 = 	 1'b0
;    6569		:	dataRd	 = 	 1'b0
;    6570		:	dataRd	 = 	 1'b0
;    6571		:	dataRd	 = 	 1'b0
;    6572		:	dataRd	 = 	 1'b0
;    6573		:	dataRd	 = 	 1'b0
;    6574		:	dataRd	 = 	 1'b0
;    6575		:	dataRd	 = 	 1'b0
;    6576		:	dataRd	 = 	 1'b0
;    6577		:	dataRd	 = 	 1'b0
;    6578		:	dataRd	 = 	 1'b0
;    6579		:	dataRd	 = 	 1'b0
;    6580		:	dataRd	 = 	 1'b0
;    6581		:	dataRd	 = 	 1'b0
;    6582		:	dataRd	 = 	 1'b0
;    6583		:	dataRd	 = 	 1'b0
;    6584		:	dataRd	 = 	 1'b0
;    6585		:	dataRd	 = 	 1'b0
;    6586		:	dataRd	 = 	 1'b0
;    6587		:	dataRd	 = 	 1'b0
;    6588		:	dataRd	 = 	 1'b0
;    6589		:	dataRd	 = 	 1'b0
;    6590		:	dataRd	 = 	 1'b0
;    6591		:	dataRd	 = 	 1'b0
;    6592		:	dataRd	 = 	 1'b0
;    6593		:	dataRd	 = 	 1'b0
;    6594		:	dataRd	 = 	 1'b0
;    6595		:	dataRd	 = 	 1'b0
;    6596		:	dataRd	 = 	 1'b0
;    6597		:	dataRd	 = 	 1'b0
;    6598		:	dataRd	 = 	 1'b0
;    6599		:	dataRd	 = 	 1'b0
;    6600		:	dataRd	 = 	 1'b0
;    6601		:	dataRd	 = 	 1'b0
;    6602		:	dataRd	 = 	 1'b0
;    6603		:	dataRd	 = 	 1'b0
;    6604		:	dataRd	 = 	 1'b0
;    6605		:	dataRd	 = 	 1'b0
;    6606		:	dataRd	 = 	 1'b0
;    6607		:	dataRd	 = 	 1'b0
;    6608		:	dataRd	 = 	 1'b0
;    6609		:	dataRd	 = 	 1'b0
;    6610		:	dataRd	 = 	 1'b0
;    6611		:	dataRd	 = 	 1'b0
;    6612		:	dataRd	 = 	 1'b0
;    6613		:	dataRd	 = 	 1'b0
;    6614		:	dataRd	 = 	 1'b0
;    6615		:	dataRd	 = 	 1'b0
;    6616		:	dataRd	 = 	 1'b0
;    6617		:	dataRd	 = 	 1'b0
;    6618		:	dataRd	 = 	 1'b0
;    6619		:	dataRd	 = 	 1'b0
;    6620		:	dataRd	 = 	 1'b0
;    6621		:	dataRd	 = 	 1'b0
;    6622		:	dataRd	 = 	 1'b0
;    6623		:	dataRd	 = 	 1'b0
;    6624		:	dataRd	 = 	 1'b0
;    6625		:	dataRd	 = 	 1'b0
;    6626		:	dataRd	 = 	 1'b0
;    6627		:	dataRd	 = 	 1'b1
;    6628		:	dataRd	 = 	 1'b0
;    6629		:	dataRd	 = 	 1'b0
;    6630		:	dataRd	 = 	 1'b0
;    6631		:	dataRd	 = 	 1'b0
;    6632		:	dataRd	 = 	 1'b0
;    6633		:	dataRd	 = 	 1'b0
;    6634		:	dataRd	 = 	 1'b0
;    6635		:	dataRd	 = 	 1'b0
;    6636		:	dataRd	 = 	 1'b0
;    6637		:	dataRd	 = 	 1'b0
;    6638		:	dataRd	 = 	 1'b0
;    6639		:	dataRd	 = 	 1'b0
;    6640		:	dataRd	 = 	 1'b0
;    6641		:	dataRd	 = 	 1'b0
;    6642		:	dataRd	 = 	 1'b0
;    6643		:	dataRd	 = 	 1'b0
;    6644		:	dataRd	 = 	 1'b0
;    6645		:	dataRd	 = 	 1'b0
;    6646		:	dataRd	 = 	 1'b0
;    6647		:	dataRd	 = 	 1'b0
;    6648		:	dataRd	 = 	 1'b0
;    6649		:	dataRd	 = 	 1'b0
;    6650		:	dataRd	 = 	 1'b0
;    6651		:	dataRd	 = 	 1'b0
;    6652		:	dataRd	 = 	 1'b0
;    6653		:	dataRd	 = 	 1'b0
;    6654		:	dataRd	 = 	 1'b0
;    6655		:	dataRd	 = 	 1'b0
;    6656		:	dataRd	 = 	 1'b0
;    6657		:	dataRd	 = 	 1'b0
;    6658		:	dataRd	 = 	 1'b0
;    6659		:	dataRd	 = 	 1'b0
;    6660		:	dataRd	 = 	 1'b0
;    6661		:	dataRd	 = 	 1'b0
;    6662		:	dataRd	 = 	 1'b0
;    6663		:	dataRd	 = 	 1'b0
;    6664		:	dataRd	 = 	 1'b0
;    6665		:	dataRd	 = 	 1'b0
;    6666		:	dataRd	 = 	 1'b0
;    6667		:	dataRd	 = 	 1'b0
;    6668		:	dataRd	 = 	 1'b0
;    6669		:	dataRd	 = 	 1'b0
;    6670		:	dataRd	 = 	 1'b0
;    6671		:	dataRd	 = 	 1'b0
;    6672		:	dataRd	 = 	 1'b0
;    6673		:	dataRd	 = 	 1'b0
;    6674		:	dataRd	 = 	 1'b0
;    6675		:	dataRd	 = 	 1'b0
;    6676		:	dataRd	 = 	 1'b0
;    6677		:	dataRd	 = 	 1'b0
;    6678		:	dataRd	 = 	 1'b0
;    6679		:	dataRd	 = 	 1'b0
;    6680		:	dataRd	 = 	 1'b0
;    6681		:	dataRd	 = 	 1'b0
;    6682		:	dataRd	 = 	 1'b0
;    6683		:	dataRd	 = 	 1'b0
;    6684		:	dataRd	 = 	 1'b0
;    6685		:	dataRd	 = 	 1'b0
;    6686		:	dataRd	 = 	 1'b0
;    6687		:	dataRd	 = 	 1'b0
;    6688		:	dataRd	 = 	 1'b0
;    6689		:	dataRd	 = 	 1'b0
;    6690		:	dataRd	 = 	 1'b0
;    6691		:	dataRd	 = 	 1'b0
;    6692		:	dataRd	 = 	 1'b0
;    6693		:	dataRd	 = 	 1'b0
;    6694		:	dataRd	 = 	 1'b1
;    6695		:	dataRd	 = 	 1'b0
;    6696		:	dataRd	 = 	 1'b0
;    6697		:	dataRd	 = 	 1'b0
;    6698		:	dataRd	 = 	 1'b0
;    6699		:	dataRd	 = 	 1'b0
;    6700		:	dataRd	 = 	 1'b0
;    6701		:	dataRd	 = 	 1'b0
;    6702		:	dataRd	 = 	 1'b0
;    6703		:	dataRd	 = 	 1'b0
;    6704		:	dataRd	 = 	 1'b0
;    6705		:	dataRd	 = 	 1'b0
;    6706		:	dataRd	 = 	 1'b0
;    6707		:	dataRd	 = 	 1'b0
;    6708		:	dataRd	 = 	 1'b0
;    6709		:	dataRd	 = 	 1'b0
;    6710		:	dataRd	 = 	 1'b0
;    6711		:	dataRd	 = 	 1'b0
;    6712		:	dataRd	 = 	 1'b0
;    6713		:	dataRd	 = 	 1'b0
;    6714		:	dataRd	 = 	 1'b0
;    6715		:	dataRd	 = 	 1'b0
;    6716		:	dataRd	 = 	 1'b0
;    6717		:	dataRd	 = 	 1'b0
;    6718		:	dataRd	 = 	 1'b0
;    6719		:	dataRd	 = 	 1'b0
;    6720		:	dataRd	 = 	 1'b0
;    6721		:	dataRd	 = 	 1'b0
;    6722		:	dataRd	 = 	 1'b0
;    6723		:	dataRd	 = 	 1'b0
;    6724		:	dataRd	 = 	 1'b0
;    6725		:	dataRd	 = 	 1'b0
;    6726		:	dataRd	 = 	 1'b0
;    6727		:	dataRd	 = 	 1'b0
;    6728		:	dataRd	 = 	 1'b0
;    6729		:	dataRd	 = 	 1'b0
;    6730		:	dataRd	 = 	 1'b0
;    6731		:	dataRd	 = 	 1'b0
;    6732		:	dataRd	 = 	 1'b0
;    6733		:	dataRd	 = 	 1'b0
;    6734		:	dataRd	 = 	 1'b0
;    6735		:	dataRd	 = 	 1'b0
;    6736		:	dataRd	 = 	 1'b0
;    6737		:	dataRd	 = 	 1'b0
;    6738		:	dataRd	 = 	 1'b0
;    6739		:	dataRd	 = 	 1'b0
;    6740		:	dataRd	 = 	 1'b0
;    6741		:	dataRd	 = 	 1'b0
;    6742		:	dataRd	 = 	 1'b0
;    6743		:	dataRd	 = 	 1'b0
;    6744		:	dataRd	 = 	 1'b0
;    6745		:	dataRd	 = 	 1'b0
;    6746		:	dataRd	 = 	 1'b0
;    6747		:	dataRd	 = 	 1'b0
;    6748		:	dataRd	 = 	 1'b0
;    6749		:	dataRd	 = 	 1'b0
;    6750		:	dataRd	 = 	 1'b0
;    6751		:	dataRd	 = 	 1'b0
;    6752		:	dataRd	 = 	 1'b0
;    6753		:	dataRd	 = 	 1'b0
;    6754		:	dataRd	 = 	 1'b0
;    6755		:	dataRd	 = 	 1'b0
;    6756		:	dataRd	 = 	 1'b0
;    6757		:	dataRd	 = 	 1'b0
;    6758		:	dataRd	 = 	 1'b0
;    6759		:	dataRd	 = 	 1'b0
;    6760		:	dataRd	 = 	 1'b0
;    6761		:	dataRd	 = 	 1'b1
;    6762		:	dataRd	 = 	 1'b0
;    6763		:	dataRd	 = 	 1'b0
;    6764		:	dataRd	 = 	 1'b0
;    6765		:	dataRd	 = 	 1'b0
;    6766		:	dataRd	 = 	 1'b0
;    6767		:	dataRd	 = 	 1'b0
;    6768		:	dataRd	 = 	 1'b0
;    6769		:	dataRd	 = 	 1'b0
;    6770		:	dataRd	 = 	 1'b0
;    6771		:	dataRd	 = 	 1'b0
;    6772		:	dataRd	 = 	 1'b0
;    6773		:	dataRd	 = 	 1'b0
;    6774		:	dataRd	 = 	 1'b0
;    6775		:	dataRd	 = 	 1'b0
;    6776		:	dataRd	 = 	 1'b0
;    6777		:	dataRd	 = 	 1'b0
;    6778		:	dataRd	 = 	 1'b0
;    6779		:	dataRd	 = 	 1'b0
;    6780		:	dataRd	 = 	 1'b0
;    6781		:	dataRd	 = 	 1'b0
;    6782		:	dataRd	 = 	 1'b0
;    6783		:	dataRd	 = 	 1'b0
;    6784		:	dataRd	 = 	 1'b0
;    6785		:	dataRd	 = 	 1'b0
;    6786		:	dataRd	 = 	 1'b0
;    6787		:	dataRd	 = 	 1'b0
;    6788		:	dataRd	 = 	 1'b0
;    6789		:	dataRd	 = 	 1'b0
;    6790		:	dataRd	 = 	 1'b0
;    6791		:	dataRd	 = 	 1'b0
;    6792		:	dataRd	 = 	 1'b0
;    6793		:	dataRd	 = 	 1'b0
;    6794		:	dataRd	 = 	 1'b0
;    6795		:	dataRd	 = 	 1'b0
;    6796		:	dataRd	 = 	 1'b0
;    6797		:	dataRd	 = 	 1'b0
;    6798		:	dataRd	 = 	 1'b0
;    6799		:	dataRd	 = 	 1'b0
;    6800		:	dataRd	 = 	 1'b0
;    6801		:	dataRd	 = 	 1'b0
;    6802		:	dataRd	 = 	 1'b0
;    6803		:	dataRd	 = 	 1'b0
;    6804		:	dataRd	 = 	 1'b0
;    6805		:	dataRd	 = 	 1'b0
;    6806		:	dataRd	 = 	 1'b0
;    6807		:	dataRd	 = 	 1'b0
;    6808		:	dataRd	 = 	 1'b0
;    6809		:	dataRd	 = 	 1'b0
;    6810		:	dataRd	 = 	 1'b0
;    6811		:	dataRd	 = 	 1'b0
;    6812		:	dataRd	 = 	 1'b0
;    6813		:	dataRd	 = 	 1'b0
;    6814		:	dataRd	 = 	 1'b0
;    6815		:	dataRd	 = 	 1'b0
;    6816		:	dataRd	 = 	 1'b0
;    6817		:	dataRd	 = 	 1'b0
;    6818		:	dataRd	 = 	 1'b0
;    6819		:	dataRd	 = 	 1'b0
;    6820		:	dataRd	 = 	 1'b0
;    6821		:	dataRd	 = 	 1'b0
;    6822		:	dataRd	 = 	 1'b0
;    6823		:	dataRd	 = 	 1'b0
;    6824		:	dataRd	 = 	 1'b0
;    6825		:	dataRd	 = 	 1'b0
;    6826		:	dataRd	 = 	 1'b0
;    6827		:	dataRd	 = 	 1'b0
;    6828		:	dataRd	 = 	 1'b0
;    6829		:	dataRd	 = 	 1'b0
;    6830		:	dataRd	 = 	 1'b0
;    6831		:	dataRd	 = 	 1'b0
;    6832		:	dataRd	 = 	 1'b0
;    6833		:	dataRd	 = 	 1'b0
;    6834		:	dataRd	 = 	 1'b0
;    6835		:	dataRd	 = 	 1'b0
;    6836		:	dataRd	 = 	 1'b0
;    6837		:	dataRd	 = 	 1'b0
;    6838		:	dataRd	 = 	 1'b0
;    6839		:	dataRd	 = 	 1'b0
;    6840		:	dataRd	 = 	 1'b0
;    6841		:	dataRd	 = 	 1'b0
;    6842		:	dataRd	 = 	 1'b0
;    6843		:	dataRd	 = 	 1'b0
;    6844		:	dataRd	 = 	 1'b0
;    6845		:	dataRd	 = 	 1'b0
;    6846		:	dataRd	 = 	 1'b0
;    6847		:	dataRd	 = 	 1'b0
;    6848		:	dataRd	 = 	 1'b0
;    6849		:	dataRd	 = 	 1'b0
;    6850		:	dataRd	 = 	 1'b0
;    6851		:	dataRd	 = 	 1'b0
;    6852		:	dataRd	 = 	 1'b0
;    6853		:	dataRd	 = 	 1'b0
;    6854		:	dataRd	 = 	 1'b0
;    6855		:	dataRd	 = 	 1'b0
;    6856		:	dataRd	 = 	 1'b0
;    6857		:	dataRd	 = 	 1'b0
;    6858		:	dataRd	 = 	 1'b0
;    6859		:	dataRd	 = 	 1'b0
;    6860		:	dataRd	 = 	 1'b0
;    6861		:	dataRd	 = 	 1'b0
;    6862		:	dataRd	 = 	 1'b0
;    6863		:	dataRd	 = 	 1'b0
;    6864		:	dataRd	 = 	 1'b0
;    6865		:	dataRd	 = 	 1'b0
;    6866		:	dataRd	 = 	 1'b0
;    6867		:	dataRd	 = 	 1'b0
;    6868		:	dataRd	 = 	 1'b0
;    6869		:	dataRd	 = 	 1'b0
;    6870		:	dataRd	 = 	 1'b0
;    6871		:	dataRd	 = 	 1'b0
;    6872		:	dataRd	 = 	 1'b0
;    6873		:	dataRd	 = 	 1'b0
;    6874		:	dataRd	 = 	 1'b0
;    6875		:	dataRd	 = 	 1'b0
;    6876		:	dataRd	 = 	 1'b0
;    6877		:	dataRd	 = 	 1'b0
;    6878		:	dataRd	 = 	 1'b0
;    6879		:	dataRd	 = 	 1'b0
;    6880		:	dataRd	 = 	 1'b0
;    6881		:	dataRd	 = 	 1'b0
;    6882		:	dataRd	 = 	 1'b0
;    6883		:	dataRd	 = 	 1'b0
;    6884		:	dataRd	 = 	 1'b0
;    6885		:	dataRd	 = 	 1'b0
;    6886		:	dataRd	 = 	 1'b0
;    6887		:	dataRd	 = 	 1'b0
;    6888		:	dataRd	 = 	 1'b1
;    6889		:	dataRd	 = 	 1'b0
;    6890		:	dataRd	 = 	 1'b0
;    6891		:	dataRd	 = 	 1'b1
;    6892		:	dataRd	 = 	 1'b0
;    6893		:	dataRd	 = 	 1'b0
;    6894		:	dataRd	 = 	 1'b1
;    6895		:	dataRd	 = 	 1'b0
;    6896		:	dataRd	 = 	 1'b0
;    6897		:	dataRd	 = 	 1'b0
;    6898		:	dataRd	 = 	 1'b0
;    6899		:	dataRd	 = 	 1'b0
;    6900		:	dataRd	 = 	 1'b0
;    6901		:	dataRd	 = 	 1'b0
;    6902		:	dataRd	 = 	 1'b0
;    6903		:	dataRd	 = 	 1'b0
;    6904		:	dataRd	 = 	 1'b0
;    6905		:	dataRd	 = 	 1'b1
;    6906		:	dataRd	 = 	 1'b0
;    6907		:	dataRd	 = 	 1'b0
;    6908		:	dataRd	 = 	 1'b0
;    6909		:	dataRd	 = 	 1'b1
;    6910		:	dataRd	 = 	 1'b1
;    6911		:	dataRd	 = 	 1'b0
;    6912		:	dataRd	 = 	 1'b0
;    6913		:	dataRd	 = 	 1'b0
;    6914		:	dataRd	 = 	 1'b0
;    6915		:	dataRd	 = 	 1'b0
;    6916		:	dataRd	 = 	 1'b0
;    6917		:	dataRd	 = 	 1'b0
;    6918		:	dataRd	 = 	 1'b1
;    6919		:	dataRd	 = 	 1'b0
;    6920		:	dataRd	 = 	 1'b0
;    6921		:	dataRd	 = 	 1'b0
;    6922		:	dataRd	 = 	 1'b0
;    6923		:	dataRd	 = 	 1'b0
;    6924		:	dataRd	 = 	 1'b0
;    6925		:	dataRd	 = 	 1'b0
;    6926		:	dataRd	 = 	 1'b0
;    6927		:	dataRd	 = 	 1'b0
;    6928		:	dataRd	 = 	 1'b1
;    6929		:	dataRd	 = 	 1'b0
;    6930		:	dataRd	 = 	 1'b0
;    6931		:	dataRd	 = 	 1'b0
;    6932		:	dataRd	 = 	 1'b0
;    6933		:	dataRd	 = 	 1'b0
;    6934		:	dataRd	 = 	 1'b1
;    6935		:	dataRd	 = 	 1'b1
;    6936		:	dataRd	 = 	 1'b1
;    6937		:	dataRd	 = 	 1'b1
;    6938		:	dataRd	 = 	 1'b1
;    6939		:	dataRd	 = 	 1'b1
;    6940		:	dataRd	 = 	 1'b1
;    6941		:	dataRd	 = 	 1'b1
;    6942		:	dataRd	 = 	 1'b0
;    6943		:	dataRd	 = 	 1'b0
;    6944		:	dataRd	 = 	 1'b0
;    6945		:	dataRd	 = 	 1'b0
;    6946		:	dataRd	 = 	 1'b0
;    6947		:	dataRd	 = 	 1'b0
;    6948		:	dataRd	 = 	 1'b0
;    6949		:	dataRd	 = 	 1'b0
;    6950		:	dataRd	 = 	 1'b0
;    6951		:	dataRd	 = 	 1'b0
;    6952		:	dataRd	 = 	 1'b0
;    6953		:	dataRd	 = 	 1'b0
;    6954		:	dataRd	 = 	 1'b0
;    6955		:	dataRd	 = 	 1'b0
;    6956		:	dataRd	 = 	 1'b0
;    6957		:	dataRd	 = 	 1'b0
;    6958		:	dataRd	 = 	 1'b0
;    6959		:	dataRd	 = 	 1'b0
;    6960		:	dataRd	 = 	 1'b0
;    6961		:	dataRd	 = 	 1'b0
;    6962		:	dataRd	 = 	 1'b0
;    6963		:	dataRd	 = 	 1'b0
;    6964		:	dataRd	 = 	 1'b0
;    6965		:	dataRd	 = 	 1'b0
;    6966		:	dataRd	 = 	 1'b0
;    6967		:	dataRd	 = 	 1'b0
;    6968		:	dataRd	 = 	 1'b0
;    6969		:	dataRd	 = 	 1'b0
;    6970		:	dataRd	 = 	 1'b0
;    6971		:	dataRd	 = 	 1'b0
;    6972		:	dataRd	 = 	 1'b0
;    6973		:	dataRd	 = 	 1'b0
;    6974		:	dataRd	 = 	 1'b0
;    6975		:	dataRd	 = 	 1'b0
;    6976		:	dataRd	 = 	 1'b0
;    6977		:	dataRd	 = 	 1'b0
;    6978		:	dataRd	 = 	 1'b1
;    6979		:	dataRd	 = 	 1'b1
;    6980		:	dataRd	 = 	 1'b0
;    6981		:	dataRd	 = 	 1'b0
;    6982		:	dataRd	 = 	 1'b0
;    6983		:	dataRd	 = 	 1'b0
;    6984		:	dataRd	 = 	 1'b0
;    6985		:	dataRd	 = 	 1'b0
;    6986		:	dataRd	 = 	 1'b0
;    6987		:	dataRd	 = 	 1'b0
;    6988		:	dataRd	 = 	 1'b0
;    6989		:	dataRd	 = 	 1'b0
;    6990		:	dataRd	 = 	 1'b0
;    6991		:	dataRd	 = 	 1'b0
;    6992		:	dataRd	 = 	 1'b1
;    6993		:	dataRd	 = 	 1'b1
;    6994		:	dataRd	 = 	 1'b1
;    6995		:	dataRd	 = 	 1'b1
;    6996		:	dataRd	 = 	 1'b1
;    6997		:	dataRd	 = 	 1'b1
;    6998		:	dataRd	 = 	 1'b1
;    6999		:	dataRd	 = 	 1'b1
;    7000		:	dataRd	 = 	 1'b0
;    7001		:	dataRd	 = 	 1'b0
;    7002		:	dataRd	 = 	 1'b0
;    7003		:	dataRd	 = 	 1'b0
;    7004		:	dataRd	 = 	 1'b0
;    7005		:	dataRd	 = 	 1'b0
;    7006		:	dataRd	 = 	 1'b0
;    7007		:	dataRd	 = 	 1'b0
;    7008		:	dataRd	 = 	 1'b0
;    7009		:	dataRd	 = 	 1'b0
;    7010		:	dataRd	 = 	 1'b0
;    7011		:	dataRd	 = 	 1'b0
;    7012		:	dataRd	 = 	 1'b0
;    7013		:	dataRd	 = 	 1'b0
;    7014		:	dataRd	 = 	 1'b0
;    7015		:	dataRd	 = 	 1'b0
;    7016		:	dataRd	 = 	 1'b0
;    7017		:	dataRd	 = 	 1'b0
;    7018		:	dataRd	 = 	 1'b0
;    7019		:	dataRd	 = 	 1'b0
;    7020		:	dataRd	 = 	 1'b0
;    7021		:	dataRd	 = 	 1'b0
;    7022		:	dataRd	 = 	 1'b0
;    7023		:	dataRd	 = 	 1'b0
;    7024		:	dataRd	 = 	 1'b0
;    7025		:	dataRd	 = 	 1'b0
;    7026		:	dataRd	 = 	 1'b0
;    7027		:	dataRd	 = 	 1'b0
;    7028		:	dataRd	 = 	 1'b0
;    7029		:	dataRd	 = 	 1'b0
;    7030		:	dataRd	 = 	 1'b1
;    7031		:	dataRd	 = 	 1'b0
;    7032		:	dataRd	 = 	 1'b0
;    7033		:	dataRd	 = 	 1'b1
;    7034		:	dataRd	 = 	 1'b0
;    7035		:	dataRd	 = 	 1'b0
;    7036		:	dataRd	 = 	 1'b0
;    7037		:	dataRd	 = 	 1'b0
;    7038		:	dataRd	 = 	 1'b1
;    7039		:	dataRd	 = 	 1'b0
;    7040		:	dataRd	 = 	 1'b0
;    7041		:	dataRd	 = 	 1'b1
;    7042		:	dataRd	 = 	 1'b0
;    7043		:	dataRd	 = 	 1'b0
;    7044		:	dataRd	 = 	 1'b1
;    7045		:	dataRd	 = 	 1'b0
;    7046		:	dataRd	 = 	 1'b0
;    7047		:	dataRd	 = 	 1'b0
;    7048		:	dataRd	 = 	 1'b0
;    7049		:	dataRd	 = 	 1'b0
;    7050		:	dataRd	 = 	 1'b1
;    7051		:	dataRd	 = 	 1'b0
;    7052		:	dataRd	 = 	 1'b0
;    7053		:	dataRd	 = 	 1'b0
;    7054		:	dataRd	 = 	 1'b0
;    7055		:	dataRd	 = 	 1'b0
;    7056		:	dataRd	 = 	 1'b1
;    7057		:	dataRd	 = 	 1'b0
;    7058		:	dataRd	 = 	 1'b0
;    7059		:	dataRd	 = 	 1'b0
;    7060		:	dataRd	 = 	 1'b0
;    7061		:	dataRd	 = 	 1'b0
;    7062		:	dataRd	 = 	 1'b1
;    7063		:	dataRd	 = 	 1'b0
;    7064		:	dataRd	 = 	 1'b0
;    7065		:	dataRd	 = 	 1'b0
;    7066		:	dataRd	 = 	 1'b0
;    7067		:	dataRd	 = 	 1'b0
;    7068		:	dataRd	 = 	 1'b0
;    7069		:	dataRd	 = 	 1'b0
;    7070		:	dataRd	 = 	 1'b1
;    7071		:	dataRd	 = 	 1'b0
;    7072		:	dataRd	 = 	 1'b0
;    7073		:	dataRd	 = 	 1'b0
;    7074		:	dataRd	 = 	 1'b0
;    7075		:	dataRd	 = 	 1'b0
;    7076		:	dataRd	 = 	 1'b0
;    7077		:	dataRd	 = 	 1'b0
;    7078		:	dataRd	 = 	 1'b0
;    7079		:	dataRd	 = 	 1'b0
;    7080		:	dataRd	 = 	 1'b0
;    7081		:	dataRd	 = 	 1'b0
;    7082		:	dataRd	 = 	 1'b0
;    7083		:	dataRd	 = 	 1'b0
;    7084		:	dataRd	 = 	 1'b0
;    7085		:	dataRd	 = 	 1'b0
;    7086		:	dataRd	 = 	 1'b0
;    7087		:	dataRd	 = 	 1'b0
;    7088		:	dataRd	 = 	 1'b0
;    7089		:	dataRd	 = 	 1'b0
;    7090		:	dataRd	 = 	 1'b0
;    7091		:	dataRd	 = 	 1'b0
;    7092		:	dataRd	 = 	 1'b0
;    7093		:	dataRd	 = 	 1'b0
;    7094		:	dataRd	 = 	 1'b0
;    7095		:	dataRd	 = 	 1'b0
;    7096		:	dataRd	 = 	 1'b1
;    7097		:	dataRd	 = 	 1'b0
;    7098		:	dataRd	 = 	 1'b0
;    7099		:	dataRd	 = 	 1'b0
;    7100		:	dataRd	 = 	 1'b0
;    7101		:	dataRd	 = 	 1'b0
;    7102		:	dataRd	 = 	 1'b1
;    7103		:	dataRd	 = 	 1'b1
;    7104		:	dataRd	 = 	 1'b1
;    7105		:	dataRd	 = 	 1'b1
;    7106		:	dataRd	 = 	 1'b1
;    7107		:	dataRd	 = 	 1'b1
;    7108		:	dataRd	 = 	 1'b1
;    7109		:	dataRd	 = 	 1'b1
;    7110		:	dataRd	 = 	 1'b0
;    7111		:	dataRd	 = 	 1'b0
;    7112		:	dataRd	 = 	 1'b0
;    7113		:	dataRd	 = 	 1'b0
;    7114		:	dataRd	 = 	 1'b0
;    7115		:	dataRd	 = 	 1'b0
;    7116		:	dataRd	 = 	 1'b0
;    7117		:	dataRd	 = 	 1'b0
;    7118		:	dataRd	 = 	 1'b0
;    7119		:	dataRd	 = 	 1'b0
;    7120		:	dataRd	 = 	 1'b0
;    7121		:	dataRd	 = 	 1'b0
;    7122		:	dataRd	 = 	 1'b0
;    7123		:	dataRd	 = 	 1'b0
;    7124		:	dataRd	 = 	 1'b0
;    7125		:	dataRd	 = 	 1'b0
;    7126		:	dataRd	 = 	 1'b0
;    7127		:	dataRd	 = 	 1'b0
;    7128		:	dataRd	 = 	 1'b0
;    7129		:	dataRd	 = 	 1'b0
;    7130		:	dataRd	 = 	 1'b0
;    7131		:	dataRd	 = 	 1'b0
;    7132		:	dataRd	 = 	 1'b0
;    7133		:	dataRd	 = 	 1'b0
;    7134		:	dataRd	 = 	 1'b0
;    7135		:	dataRd	 = 	 1'b0
;    7136		:	dataRd	 = 	 1'b0
;    7137		:	dataRd	 = 	 1'b0
;    7138		:	dataRd	 = 	 1'b0
;    7139		:	dataRd	 = 	 1'b0
;    7140		:	dataRd	 = 	 1'b0
;    7141		:	dataRd	 = 	 1'b0
;    7142		:	dataRd	 = 	 1'b0
;    7143		:	dataRd	 = 	 1'b0
;    7144		:	dataRd	 = 	 1'b1
;    7145		:	dataRd	 = 	 1'b0
;    7146		:	dataRd	 = 	 1'b0
;    7147		:	dataRd	 = 	 1'b0
;    7148		:	dataRd	 = 	 1'b0
;    7149		:	dataRd	 = 	 1'b0
;    7150		:	dataRd	 = 	 1'b0
;    7151		:	dataRd	 = 	 1'b0
;    7152		:	dataRd	 = 	 1'b1
;    7153		:	dataRd	 = 	 1'b0
;    7154		:	dataRd	 = 	 1'b0
;    7155		:	dataRd	 = 	 1'b0
;    7156		:	dataRd	 = 	 1'b0
;    7157		:	dataRd	 = 	 1'b0
;    7158		:	dataRd	 = 	 1'b0
;    7159		:	dataRd	 = 	 1'b0
;    7160		:	dataRd	 = 	 1'b0
;    7161		:	dataRd	 = 	 1'b0
;    7162		:	dataRd	 = 	 1'b0
;    7163		:	dataRd	 = 	 1'b0
;    7164		:	dataRd	 = 	 1'b0
;    7165		:	dataRd	 = 	 1'b0
;    7166		:	dataRd	 = 	 1'b0
;    7167		:	dataRd	 = 	 1'b0
;    7168		:	dataRd	 = 	 1'b0
;    7169		:	dataRd	 = 	 1'b0
;    7170		:	dataRd	 = 	 1'b1
;    7171		:	dataRd	 = 	 1'b0
;    7172		:	dataRd	 = 	 1'b0
;    7173		:	dataRd	 = 	 1'b1
;    7174		:	dataRd	 = 	 1'b0
;    7175		:	dataRd	 = 	 1'b0
;    7176		:	dataRd	 = 	 1'b1
;    7177		:	dataRd	 = 	 1'b0
;    7178		:	dataRd	 = 	 1'b0
;    7179		:	dataRd	 = 	 1'b0
;    7180		:	dataRd	 = 	 1'b0
;    7181		:	dataRd	 = 	 1'b0
;    7182		:	dataRd	 = 	 1'b0
;    7183		:	dataRd	 = 	 1'b0
;    7184		:	dataRd	 = 	 1'b1
;    7185		:	dataRd	 = 	 1'b1
;    7186		:	dataRd	 = 	 1'b1
;    7187		:	dataRd	 = 	 1'b1
;    7188		:	dataRd	 = 	 1'b1
;    7189		:	dataRd	 = 	 1'b1
;    7190		:	dataRd	 = 	 1'b1
;    7191		:	dataRd	 = 	 1'b1
;    7192		:	dataRd	 = 	 1'b0
;    7193		:	dataRd	 = 	 1'b0
;    7194		:	dataRd	 = 	 1'b0
;    7195		:	dataRd	 = 	 1'b0
;    7196		:	dataRd	 = 	 1'b0
;    7197		:	dataRd	 = 	 1'b0
;    7198		:	dataRd	 = 	 1'b0
;    7199		:	dataRd	 = 	 1'b0
;    7200		:	dataRd	 = 	 1'b0
;    7201		:	dataRd	 = 	 1'b0
;    7202		:	dataRd	 = 	 1'b0
;    7203		:	dataRd	 = 	 1'b0
;    7204		:	dataRd	 = 	 1'b0
;    7205		:	dataRd	 = 	 1'b0
;    7206		:	dataRd	 = 	 1'b0
;    7207		:	dataRd	 = 	 1'b0
;    7208		:	dataRd	 = 	 1'b0
;    7209		:	dataRd	 = 	 1'b0
;    7210		:	dataRd	 = 	 1'b0
;    7211		:	dataRd	 = 	 1'b0
;    7212		:	dataRd	 = 	 1'b0
;    7213		:	dataRd	 = 	 1'b0
;    7214		:	dataRd	 = 	 1'b0
;    7215		:	dataRd	 = 	 1'b0
;    7216		:	dataRd	 = 	 1'b0
;    7217		:	dataRd	 = 	 1'b0
;    7218		:	dataRd	 = 	 1'b0
;    7219		:	dataRd	 = 	 1'b0
;    7220		:	dataRd	 = 	 1'b0
;    7221		:	dataRd	 = 	 1'b0
;    7222		:	dataRd	 = 	 1'b0
;    7223		:	dataRd	 = 	 1'b0
;    7224		:	dataRd	 = 	 1'b0
;    7225		:	dataRd	 = 	 1'b0
;    7226		:	dataRd	 = 	 1'b0
;    7227		:	dataRd	 = 	 1'b0
;    7228		:	dataRd	 = 	 1'b0
;    7229		:	dataRd	 = 	 1'b0
;    7230		:	dataRd	 = 	 1'b0
;    7231		:	dataRd	 = 	 1'b0
;    7232		:	dataRd	 = 	 1'b0
;    7233		:	dataRd	 = 	 1'b0
;    7234		:	dataRd	 = 	 1'b1
;    7235		:	dataRd	 = 	 1'b0
;    7236		:	dataRd	 = 	 1'b0
;    7237		:	dataRd	 = 	 1'b0
;    7238		:	dataRd	 = 	 1'b0
;    7239		:	dataRd	 = 	 1'b0
;    7240		:	dataRd	 = 	 1'b0
;    7241		:	dataRd	 = 	 1'b0
;    7242		:	dataRd	 = 	 1'b0
;    7243		:	dataRd	 = 	 1'b0
;    7244		:	dataRd	 = 	 1'b0
;    7245		:	dataRd	 = 	 1'b0
;    7246		:	dataRd	 = 	 1'b0
;    7247		:	dataRd	 = 	 1'b0
;    7248		:	dataRd	 = 	 1'b1
;    7249		:	dataRd	 = 	 1'b0
;    7250		:	dataRd	 = 	 1'b0
;    7251		:	dataRd	 = 	 1'b0
;    7252		:	dataRd	 = 	 1'b0
;    7253		:	dataRd	 = 	 1'b0
;    7254		:	dataRd	 = 	 1'b1
;    7255		:	dataRd	 = 	 1'b1
;    7256		:	dataRd	 = 	 1'b1
;    7257		:	dataRd	 = 	 1'b1
;    7258		:	dataRd	 = 	 1'b1
;    7259		:	dataRd	 = 	 1'b1
;    7260		:	dataRd	 = 	 1'b1
;    7261		:	dataRd	 = 	 1'b1
;    7262		:	dataRd	 = 	 1'b1
;    7263		:	dataRd	 = 	 1'b1
;    7264		:	dataRd	 = 	 1'b1
;    7265		:	dataRd	 = 	 1'b1
;    7266		:	dataRd	 = 	 1'b1
;    7267		:	dataRd	 = 	 1'b1
;    7268		:	dataRd	 = 	 1'b1
;    7269		:	dataRd	 = 	 1'b1
;    7270		:	dataRd	 = 	 1'b1
;    7271		:	dataRd	 = 	 1'b1
;    7272		:	dataRd	 = 	 1'b1
;    7273		:	dataRd	 = 	 1'b1
;    7274		:	dataRd	 = 	 1'b1
;    7275		:	dataRd	 = 	 1'b0
;    7276		:	dataRd	 = 	 1'b1
;    7277		:	dataRd	 = 	 1'b1
;    7278		:	dataRd	 = 	 1'b1
;    7279		:	dataRd	 = 	 1'b1
;    7280		:	dataRd	 = 	 1'b1
;    7281		:	dataRd	 = 	 1'b1
;    7282		:	dataRd	 = 	 1'b1
;    7283		:	dataRd	 = 	 1'b1
;    7284		:	dataRd	 = 	 1'b1
;    7285		:	dataRd	 = 	 1'b1
;	 default	:	dataRd		=	1'b0;
	endcase

end

endmodule