//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][14]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Jul  6 16:45:16 2023
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for sb_0__14_ -----
module sb_0__14_(pReset,
                 prog_clk,
                 chanx_right_in,
                 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
                 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_,
                 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
                 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
                 chany_bottom_in,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_,
                 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                 ccff_head,
                 chanx_right_out,
                 chany_bottom_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:49] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:49] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:49] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:49] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_2level_tapbuf_size2_0_sram;
wire [0:1] mux_2level_tapbuf_size2_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_10_sram;
wire [0:1] mux_2level_tapbuf_size2_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_11_sram;
wire [0:1] mux_2level_tapbuf_size2_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_12_sram;
wire [0:1] mux_2level_tapbuf_size2_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_13_sram;
wire [0:1] mux_2level_tapbuf_size2_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_14_sram;
wire [0:1] mux_2level_tapbuf_size2_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_15_sram;
wire [0:1] mux_2level_tapbuf_size2_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_16_sram;
wire [0:1] mux_2level_tapbuf_size2_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_17_sram;
wire [0:1] mux_2level_tapbuf_size2_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_18_sram;
wire [0:1] mux_2level_tapbuf_size2_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_19_sram;
wire [0:1] mux_2level_tapbuf_size2_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_1_sram;
wire [0:1] mux_2level_tapbuf_size2_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_20_sram;
wire [0:1] mux_2level_tapbuf_size2_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_21_sram;
wire [0:1] mux_2level_tapbuf_size2_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_22_sram;
wire [0:1] mux_2level_tapbuf_size2_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_23_sram;
wire [0:1] mux_2level_tapbuf_size2_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_24_sram;
wire [0:1] mux_2level_tapbuf_size2_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_25_sram;
wire [0:1] mux_2level_tapbuf_size2_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_26_sram;
wire [0:1] mux_2level_tapbuf_size2_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_27_sram;
wire [0:1] mux_2level_tapbuf_size2_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_28_sram;
wire [0:1] mux_2level_tapbuf_size2_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_29_sram;
wire [0:1] mux_2level_tapbuf_size2_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_2_sram;
wire [0:1] mux_2level_tapbuf_size2_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_30_sram;
wire [0:1] mux_2level_tapbuf_size2_30_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_31_sram;
wire [0:1] mux_2level_tapbuf_size2_31_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_32_sram;
wire [0:1] mux_2level_tapbuf_size2_32_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_33_sram;
wire [0:1] mux_2level_tapbuf_size2_33_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_34_sram;
wire [0:1] mux_2level_tapbuf_size2_34_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_35_sram;
wire [0:1] mux_2level_tapbuf_size2_35_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_36_sram;
wire [0:1] mux_2level_tapbuf_size2_36_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_37_sram;
wire [0:1] mux_2level_tapbuf_size2_37_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_38_sram;
wire [0:1] mux_2level_tapbuf_size2_38_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_39_sram;
wire [0:1] mux_2level_tapbuf_size2_39_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_3_sram;
wire [0:1] mux_2level_tapbuf_size2_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_40_sram;
wire [0:1] mux_2level_tapbuf_size2_40_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_41_sram;
wire [0:1] mux_2level_tapbuf_size2_41_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_42_sram;
wire [0:1] mux_2level_tapbuf_size2_42_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_43_sram;
wire [0:1] mux_2level_tapbuf_size2_43_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_44_sram;
wire [0:1] mux_2level_tapbuf_size2_44_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_45_sram;
wire [0:1] mux_2level_tapbuf_size2_45_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_46_sram;
wire [0:1] mux_2level_tapbuf_size2_46_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_47_sram;
wire [0:1] mux_2level_tapbuf_size2_47_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_48_sram;
wire [0:1] mux_2level_tapbuf_size2_48_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_49_sram;
wire [0:1] mux_2level_tapbuf_size2_49_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_4_sram;
wire [0:1] mux_2level_tapbuf_size2_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_50_sram;
wire [0:1] mux_2level_tapbuf_size2_50_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_51_sram;
wire [0:1] mux_2level_tapbuf_size2_51_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_52_sram;
wire [0:1] mux_2level_tapbuf_size2_52_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_53_sram;
wire [0:1] mux_2level_tapbuf_size2_53_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_54_sram;
wire [0:1] mux_2level_tapbuf_size2_54_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_55_sram;
wire [0:1] mux_2level_tapbuf_size2_55_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_56_sram;
wire [0:1] mux_2level_tapbuf_size2_56_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_57_sram;
wire [0:1] mux_2level_tapbuf_size2_57_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_58_sram;
wire [0:1] mux_2level_tapbuf_size2_58_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_59_sram;
wire [0:1] mux_2level_tapbuf_size2_59_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_5_sram;
wire [0:1] mux_2level_tapbuf_size2_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_60_sram;
wire [0:1] mux_2level_tapbuf_size2_60_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_61_sram;
wire [0:1] mux_2level_tapbuf_size2_61_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_62_sram;
wire [0:1] mux_2level_tapbuf_size2_62_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_63_sram;
wire [0:1] mux_2level_tapbuf_size2_63_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_64_sram;
wire [0:1] mux_2level_tapbuf_size2_64_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_65_sram;
wire [0:1] mux_2level_tapbuf_size2_65_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_66_sram;
wire [0:1] mux_2level_tapbuf_size2_66_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_67_sram;
wire [0:1] mux_2level_tapbuf_size2_67_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_68_sram;
wire [0:1] mux_2level_tapbuf_size2_68_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_69_sram;
wire [0:1] mux_2level_tapbuf_size2_69_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_6_sram;
wire [0:1] mux_2level_tapbuf_size2_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_7_sram;
wire [0:1] mux_2level_tapbuf_size2_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_8_sram;
wire [0:1] mux_2level_tapbuf_size2_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size2_9_sram;
wire [0:1] mux_2level_tapbuf_size2_9_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_0_sram;
wire [0:1] mux_2level_tapbuf_size3_0_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_10_sram;
wire [0:1] mux_2level_tapbuf_size3_10_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_11_sram;
wire [0:1] mux_2level_tapbuf_size3_11_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_12_sram;
wire [0:1] mux_2level_tapbuf_size3_12_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_13_sram;
wire [0:1] mux_2level_tapbuf_size3_13_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_14_sram;
wire [0:1] mux_2level_tapbuf_size3_14_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_15_sram;
wire [0:1] mux_2level_tapbuf_size3_15_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_16_sram;
wire [0:1] mux_2level_tapbuf_size3_16_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_17_sram;
wire [0:1] mux_2level_tapbuf_size3_17_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_18_sram;
wire [0:1] mux_2level_tapbuf_size3_18_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_19_sram;
wire [0:1] mux_2level_tapbuf_size3_19_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_1_sram;
wire [0:1] mux_2level_tapbuf_size3_1_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_20_sram;
wire [0:1] mux_2level_tapbuf_size3_20_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_21_sram;
wire [0:1] mux_2level_tapbuf_size3_21_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_22_sram;
wire [0:1] mux_2level_tapbuf_size3_22_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_23_sram;
wire [0:1] mux_2level_tapbuf_size3_23_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_24_sram;
wire [0:1] mux_2level_tapbuf_size3_24_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_25_sram;
wire [0:1] mux_2level_tapbuf_size3_25_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_26_sram;
wire [0:1] mux_2level_tapbuf_size3_26_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_27_sram;
wire [0:1] mux_2level_tapbuf_size3_27_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_28_sram;
wire [0:1] mux_2level_tapbuf_size3_28_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_29_sram;
wire [0:1] mux_2level_tapbuf_size3_29_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_2_sram;
wire [0:1] mux_2level_tapbuf_size3_2_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_3_sram;
wire [0:1] mux_2level_tapbuf_size3_3_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_4_sram;
wire [0:1] mux_2level_tapbuf_size3_4_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_5_sram;
wire [0:1] mux_2level_tapbuf_size3_5_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_6_sram;
wire [0:1] mux_2level_tapbuf_size3_6_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_7_sram;
wire [0:1] mux_2level_tapbuf_size3_7_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_8_sram;
wire [0:1] mux_2level_tapbuf_size3_8_sram_inv;
wire [0:1] mux_2level_tapbuf_size3_9_sram;
wire [0:1] mux_2level_tapbuf_size3_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_2level_tapbuf_size3 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[48]}),
		.sram(mux_2level_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_2level_tapbuf_size3 mux_right_track_2 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[47]}),
		.sram(mux_2level_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_2level_tapbuf_size3 mux_right_track_4 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[46]}),
		.sram(mux_2level_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_2level_tapbuf_size3 mux_right_track_20 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[38]}),
		.sram(mux_2level_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_2level_tapbuf_size3 mux_right_track_22 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[37]}),
		.sram(mux_2level_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_2level_tapbuf_size3 mux_right_track_24 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[36]}),
		.sram(mux_2level_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_2level_tapbuf_size3 mux_right_track_40 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[28]}),
		.sram(mux_2level_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_2level_tapbuf_size3 mux_right_track_42 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[27]}),
		.sram(mux_2level_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_2level_tapbuf_size3 mux_right_track_44 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[26]}),
		.sram(mux_2level_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_2level_tapbuf_size3 mux_right_track_60 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[18]}),
		.sram(mux_2level_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_2level_tapbuf_size3 mux_right_track_62 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[17]}),
		.sram(mux_2level_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_2level_tapbuf_size3 mux_right_track_64 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[16]}),
		.sram(mux_2level_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_2level_tapbuf_size3 mux_right_track_80 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_, chany_bottom_in[8]}),
		.sram(mux_2level_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_2level_tapbuf_size3 mux_right_track_82 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, chany_bottom_in[7]}),
		.sram(mux_2level_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_2level_tapbuf_size3 mux_right_track_84 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, chany_bottom_in[6]}),
		.sram(mux_2level_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_2level_tapbuf_size3 mux_bottom_track_1 (
		.in({chanx_right_in[48], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_bottom_out[0]));

	mux_2level_tapbuf_size3 mux_bottom_track_3 (
		.in({chanx_right_in[47], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_bottom_out[1]));

	mux_2level_tapbuf_size3 mux_bottom_track_5 (
		.in({chanx_right_in[46], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_bottom_out[2]));

	mux_2level_tapbuf_size3 mux_bottom_track_21 (
		.in({chanx_right_in[38], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	mux_2level_tapbuf_size3 mux_bottom_track_23 (
		.in({chanx_right_in[37], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	mux_2level_tapbuf_size3 mux_bottom_track_25 (
		.in({chanx_right_in[36], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	mux_2level_tapbuf_size3 mux_bottom_track_41 (
		.in({chanx_right_in[28], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_bottom_out[20]));

	mux_2level_tapbuf_size3 mux_bottom_track_43 (
		.in({chanx_right_in[27], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_bottom_out[21]));

	mux_2level_tapbuf_size3 mux_bottom_track_45 (
		.in({chanx_right_in[26], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_bottom_out[22]));

	mux_2level_tapbuf_size3 mux_bottom_track_61 (
		.in({chanx_right_in[18], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_bottom_out[30]));

	mux_2level_tapbuf_size3 mux_bottom_track_63 (
		.in({chanx_right_in[17], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_bottom_out[31]));

	mux_2level_tapbuf_size3 mux_bottom_track_65 (
		.in({chanx_right_in[16], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	mux_2level_tapbuf_size3 mux_bottom_track_81 (
		.in({chanx_right_in[8], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	mux_2level_tapbuf_size3 mux_bottom_track_83 (
		.in({chanx_right_in[7], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	mux_2level_tapbuf_size3 mux_bottom_track_85 (
		.in({chanx_right_in[6], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	mux_2level_tapbuf_size3_mem mem_right_track_0 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_0_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_2 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_1_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_4 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_2_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_20 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_3_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_22 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_4_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_24 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_5_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_40 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_6_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_42 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_7_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_44 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_8_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_60 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_9_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_62 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_10_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_64 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_11_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_80 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_12_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_82 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_13_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_right_track_84 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_14_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_1 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_15_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_3 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_16_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_5 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_17_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_21 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_18_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_23 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_19_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_25 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_20_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_41 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_21_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_43 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_22_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_45 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_23_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_61 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_24_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_63 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_25_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_65 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_26_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_81 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_27_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_83 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_28_sram_inv[0:1]));

	mux_2level_tapbuf_size3_mem mem_bottom_track_85 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size3_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2 mux_right_track_6 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[45]}),
		.sram(mux_2level_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_2level_tapbuf_size2 mux_right_track_8 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[44]}),
		.sram(mux_2level_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_2level_tapbuf_size2 mux_right_track_10 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[43]}),
		.sram(mux_2level_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_2level_tapbuf_size2 mux_right_track_12 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[42]}),
		.sram(mux_2level_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_2level_tapbuf_size2 mux_right_track_14 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[41]}),
		.sram(mux_2level_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_2level_tapbuf_size2 mux_right_track_16 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[40]}),
		.sram(mux_2level_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_2level_tapbuf_size2 mux_right_track_18 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[39]}),
		.sram(mux_2level_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_2level_tapbuf_size2 mux_right_track_26 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[35]}),
		.sram(mux_2level_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_2level_tapbuf_size2 mux_right_track_28 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[34]}),
		.sram(mux_2level_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_2level_tapbuf_size2 mux_right_track_30 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[33]}),
		.sram(mux_2level_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_9_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_2level_tapbuf_size2 mux_right_track_32 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[32]}),
		.sram(mux_2level_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_10_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_2level_tapbuf_size2 mux_right_track_34 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[31]}),
		.sram(mux_2level_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_11_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_2level_tapbuf_size2 mux_right_track_36 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[30]}),
		.sram(mux_2level_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_12_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_2level_tapbuf_size2 mux_right_track_38 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[29]}),
		.sram(mux_2level_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_13_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_2level_tapbuf_size2 mux_right_track_46 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[25]}),
		.sram(mux_2level_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_14_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_2level_tapbuf_size2 mux_right_track_48 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[24]}),
		.sram(mux_2level_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_15_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_2level_tapbuf_size2 mux_right_track_50 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[23]}),
		.sram(mux_2level_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_16_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_2level_tapbuf_size2 mux_right_track_52 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[22]}),
		.sram(mux_2level_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_17_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_2level_tapbuf_size2 mux_right_track_54 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[21]}),
		.sram(mux_2level_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_18_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_2level_tapbuf_size2 mux_right_track_56 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[20]}),
		.sram(mux_2level_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_19_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_2level_tapbuf_size2 mux_right_track_58 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[19]}),
		.sram(mux_2level_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_20_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_2level_tapbuf_size2 mux_right_track_66 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[15]}),
		.sram(mux_2level_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_21_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_2level_tapbuf_size2 mux_right_track_68 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[14]}),
		.sram(mux_2level_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_22_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_2level_tapbuf_size2 mux_right_track_70 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[13]}),
		.sram(mux_2level_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_23_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_2level_tapbuf_size2 mux_right_track_72 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[12]}),
		.sram(mux_2level_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_24_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_2level_tapbuf_size2 mux_right_track_74 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[11]}),
		.sram(mux_2level_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_25_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_2level_tapbuf_size2 mux_right_track_76 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[10]}),
		.sram(mux_2level_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_26_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_2level_tapbuf_size2 mux_right_track_78 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[9]}),
		.sram(mux_2level_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_27_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_2level_tapbuf_size2 mux_right_track_86 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[5]}),
		.sram(mux_2level_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_28_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_2level_tapbuf_size2 mux_right_track_88 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[4]}),
		.sram(mux_2level_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_29_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_2level_tapbuf_size2 mux_right_track_90 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[3]}),
		.sram(mux_2level_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_30_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_2level_tapbuf_size2 mux_right_track_92 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[2]}),
		.sram(mux_2level_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_31_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_2level_tapbuf_size2 mux_right_track_94 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[1]}),
		.sram(mux_2level_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_32_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_2level_tapbuf_size2 mux_right_track_96 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[0]}),
		.sram(mux_2level_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_33_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_2level_tapbuf_size2 mux_right_track_98 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_, chany_bottom_in[49]}),
		.sram(mux_2level_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_34_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_2level_tapbuf_size2 mux_bottom_track_7 (
		.in({chanx_right_in[45], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_35_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	mux_2level_tapbuf_size2 mux_bottom_track_9 (
		.in({chanx_right_in[44], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_36_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	mux_2level_tapbuf_size2 mux_bottom_track_11 (
		.in({chanx_right_in[43], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_37_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	mux_2level_tapbuf_size2 mux_bottom_track_13 (
		.in({chanx_right_in[42], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_38_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	mux_2level_tapbuf_size2 mux_bottom_track_15 (
		.in({chanx_right_in[41], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_39_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	mux_2level_tapbuf_size2 mux_bottom_track_17 (
		.in({chanx_right_in[40], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_40_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	mux_2level_tapbuf_size2 mux_bottom_track_19 (
		.in({chanx_right_in[39], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_41_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	mux_2level_tapbuf_size2 mux_bottom_track_27 (
		.in({chanx_right_in[35], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_42_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	mux_2level_tapbuf_size2 mux_bottom_track_29 (
		.in({chanx_right_in[34], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_43_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	mux_2level_tapbuf_size2 mux_bottom_track_31 (
		.in({chanx_right_in[33], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_44_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	mux_2level_tapbuf_size2 mux_bottom_track_33 (
		.in({chanx_right_in[32], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_45_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_2level_tapbuf_size2 mux_bottom_track_35 (
		.in({chanx_right_in[31], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_46_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_2level_tapbuf_size2 mux_bottom_track_37 (
		.in({chanx_right_in[30], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_47_sram_inv[0:1]),
		.out(chany_bottom_out[18]));

	mux_2level_tapbuf_size2 mux_bottom_track_39 (
		.in({chanx_right_in[29], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_48_sram_inv[0:1]),
		.out(chany_bottom_out[19]));

	mux_2level_tapbuf_size2 mux_bottom_track_47 (
		.in({chanx_right_in[25], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_49_sram_inv[0:1]),
		.out(chany_bottom_out[23]));

	mux_2level_tapbuf_size2 mux_bottom_track_49 (
		.in({chanx_right_in[24], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_50_sram_inv[0:1]),
		.out(chany_bottom_out[24]));

	mux_2level_tapbuf_size2 mux_bottom_track_51 (
		.in({chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_51_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	mux_2level_tapbuf_size2 mux_bottom_track_53 (
		.in({chanx_right_in[22], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_52_sram_inv[0:1]),
		.out(chany_bottom_out[26]));

	mux_2level_tapbuf_size2 mux_bottom_track_55 (
		.in({chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_53_sram_inv[0:1]),
		.out(chany_bottom_out[27]));

	mux_2level_tapbuf_size2 mux_bottom_track_57 (
		.in({chanx_right_in[20], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_54_sram_inv[0:1]),
		.out(chany_bottom_out[28]));

	mux_2level_tapbuf_size2 mux_bottom_track_59 (
		.in({chanx_right_in[19], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_55_sram_inv[0:1]),
		.out(chany_bottom_out[29]));

	mux_2level_tapbuf_size2 mux_bottom_track_67 (
		.in({chanx_right_in[15], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_56_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	mux_2level_tapbuf_size2 mux_bottom_track_69 (
		.in({chanx_right_in[14], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_57_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	mux_2level_tapbuf_size2 mux_bottom_track_71 (
		.in({chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_58_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	mux_2level_tapbuf_size2 mux_bottom_track_73 (
		.in({chanx_right_in[12], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_59_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	mux_2level_tapbuf_size2 mux_bottom_track_75 (
		.in({chanx_right_in[11], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_60_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	mux_2level_tapbuf_size2 mux_bottom_track_77 (
		.in({chanx_right_in[10], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_61_sram_inv[0:1]),
		.out(chany_bottom_out[38]));

	mux_2level_tapbuf_size2 mux_bottom_track_79 (
		.in({chanx_right_in[9], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_62_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	mux_2level_tapbuf_size2 mux_bottom_track_87 (
		.in({chanx_right_in[5], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(mux_2level_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_63_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	mux_2level_tapbuf_size2 mux_bottom_track_89 (
		.in({chanx_right_in[4], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(mux_2level_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_64_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	mux_2level_tapbuf_size2 mux_bottom_track_91 (
		.in({chanx_right_in[3], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_65_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	mux_2level_tapbuf_size2 mux_bottom_track_93 (
		.in({chanx_right_in[2], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_66_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	mux_2level_tapbuf_size2 mux_bottom_track_95 (
		.in({chanx_right_in[1], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_67_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	mux_2level_tapbuf_size2 mux_bottom_track_97 (
		.in({chanx_right_in[0], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_68_sram_inv[0:1]),
		.out(chany_bottom_out[48]));

	mux_2level_tapbuf_size2 mux_bottom_track_99 (
		.in({chanx_right_in[49], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_2level_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_2level_tapbuf_size2_69_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	mux_2level_tapbuf_size2_mem mem_right_track_6 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_0_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_8 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_1_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_10 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_2_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_12 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_3_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_14 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_4_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_16 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_5_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_18 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_6_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_26 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_7_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_28 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_8_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_30 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_9_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_32 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_10_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_34 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_11_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_36 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_12_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_38 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_13_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_46 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_14_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_48 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_15_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_50 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_16_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_52 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_17_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_54 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_18_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_56 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_19_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_58 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_20_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_66 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_21_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_68 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_22_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_70 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_23_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_72 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_24_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_74 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_25_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_76 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_26_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_78 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_27_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_86 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_28_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_88 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_29_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_90 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_30_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_92 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_31_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_94 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_32_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_96 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_33_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_right_track_98 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_34_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_7 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_35_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_9 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_36_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_11 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_37_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_13 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_38_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_15 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_39_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_17 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_40_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_19 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_41_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_27 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_42_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_29 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_43_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_31 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_44_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_33 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_45_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_35 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_46_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_37 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_47_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_39 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_48_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_47 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_49_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_49 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_50_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_51 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_51_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_53 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_52_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_55 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_53_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_57 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_54_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_59 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_55_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_67 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_56_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_69 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_57_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_71 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_58_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_73 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_59_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_75 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_60_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_77 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_61_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_79 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_62_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_87 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_63_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_89 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_64_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_91 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_65_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_93 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_66_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_95 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_67_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_97 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_68_sram_inv[0:1]));

	mux_2level_tapbuf_size2_mem mem_bottom_track_99 (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.ccff_head(mux_2level_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_2level_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_2level_tapbuf_size2_69_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__14_ -----

//----- Default net type -----
`default_nettype none



